
module c5315 ( N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, 
        N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, 
        N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
        N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
        N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, 
        N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, 
        N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, 
        N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
        N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, 
        N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, 
        N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, 
        N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, 
        N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
        N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, 
        N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, 
        N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, 
        N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, 
        N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, 
        N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, 
        N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, 
        N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, 
        N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, 
        N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, 
        N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, 
        N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, 
        N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, 
        N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128 );
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37,
         N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79,
         N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106,
         N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136,
         N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164,
         N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197,
         N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234,
         N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273,
         N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
         N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358,
         N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422,
         N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545,
         N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583,
         N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610,
         N613, N616, N619, N625, N631;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060,
         N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
         N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737,
         N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716,
         N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449,
         N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476,
         N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520,
         N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
         N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754,
         N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
         N8124, N8127, N8128;
  wire   N0, N6927, n1161, N1137, N1141, n485, n487, n489, n491, n493, n495,
         n497, n499, N6643, n501, N4278, n503, n504, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, N6926,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, N2527, N709, N2309, N6648;
  assign N1972 = N0;
  assign N6925 = N6927;
  assign N1143 = N1137;
  assign N1142 = N1137;
  assign N2584 = N1141;
  assign N6646 = N6643;
  assign N4275 = N4278;
  assign N6924 = N6926;
  assign N3604 = N2527;
  assign N2142 = N709;
  assign N3360 = N2309;
  assign N3359 = N2309;
  assign N3358 = N2309;
  assign N3357 = N2309;
  assign N6641 = N6648;

  HS65_LH_IVX22 U543 ( .A(n1122), .Z(N7699) );
  HS65_LH_IVX27 U544 ( .A(n497), .Z(N4272) );
  HS65_LL_IVX13 U545 ( .A(n493), .Z(N4737) );
  HS65_LH_BFX22 U546 ( .A(n988), .Z(N5240) );
  HS65_LH_AO222X4 U547 ( .A(n1113), .B(n1040), .C(n1011), .D(N117), .E(n1042), 
        .F(n699), .Z(n700) );
  HS65_LH_IVX4 U548 ( .A(N7472), .Z(n1139) );
  HS65_LH_OAI21X2 U549 ( .A(n1117), .B(n1116), .C(n1115), .Z(n1118) );
  HS65_LH_OAI12X2 U550 ( .A(n895), .B(n1049), .C(n894), .Z(n897) );
  HS65_LH_IVX9 U551 ( .A(n1095), .Z(n485) );
  HS65_LH_IVX35 U552 ( .A(n495), .Z(N2387) );
  HS65_LH_BFX49 U553 ( .A(N592), .Z(N1066) );
  HS65_LL_AO222X4 U554 ( .A(n1108), .B(n1040), .C(n1011), .D(N122), .E(n1042), 
        .F(n898), .Z(n1078) );
  HS65_LH_BFX9 U555 ( .A(n1094), .Z(n1095) );
  HS65_LH_NAND2AX7 U556 ( .A(n665), .B(n664), .Z(n1079) );
  HS65_LH_NAND2AX7 U557 ( .A(n783), .B(n782), .Z(n1114) );
  HS65_LL_NOR2X6 U558 ( .A(N616), .B(n725), .Z(n1128) );
  HS65_LL_AND2X18 U559 ( .A(N552), .B(N562), .Z(N1140) );
  HS65_LH_OAI12X18 U560 ( .A(n1002), .B(n1001), .C(n1000), .Z(n1122) );
  HS65_LH_AND2X4 U561 ( .A(N574), .B(n645), .Z(n1130) );
  HS65_LH_AND2X4 U562 ( .A(N613), .B(N616), .Z(n711) );
  HS65_LH_AND2X4 U563 ( .A(N580), .B(n668), .Z(n1134) );
  HS65_LH_NOR2X6 U564 ( .A(N574), .B(n644), .Z(n1133) );
  HS65_LH_BFX9 U565 ( .A(N549), .Z(n695) );
  HS65_LL_BFX27 U566 ( .A(N141), .Z(N709) );
  HS65_LL_AOI21X2 U567 ( .A(n992), .B(n915), .C(n738), .Z(n739) );
  HS65_LH_MUXI41X2 U568 ( .D0(N596), .D1(n1007), .D2(N595), .D3(n1006), .S0(
        N400), .S1(N265), .Z(n1109) );
  HS65_LH_AND2X4 U569 ( .A(N610), .B(N607), .Z(n1029) );
  HS65_LH_IVX9 U570 ( .A(n1040), .Z(n506) );
  HS65_LH_IVX9 U571 ( .A(n1042), .Z(n1037) );
  HS65_LH_IVX9 U572 ( .A(N2139), .Z(n1083) );
  HS65_LH_MUXI21X2 U573 ( .D0(N597), .D1(N598), .S0(N210), .Z(n727) );
  HS65_LL_OAI12X3 U574 ( .A(n570), .B(n569), .C(n568), .Z(n599) );
  HS65_LL_NOR2X13 U575 ( .A(N625), .B(n874), .Z(n1042) );
  HS65_LL_NOR2X6 U576 ( .A(N619), .B(n618), .Z(n1011) );
  HS65_LL_NOR2X6 U577 ( .A(N625), .B(N619), .Z(n1040) );
  HS65_LH_MUXI41X2 U578 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(N351), .S1(N534), .Z(n614) );
  HS65_LH_MUXI41X2 U579 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(N341), .S1(N523), .Z(n603) );
  HS65_LL_XOR2X4 U580 ( .A(n793), .B(n792), .Z(n794) );
  HS65_LL_XOR3X9 U581 ( .A(n549), .B(n716), .C(n582), .Z(n563) );
  HS65_LH_IVX9 U582 ( .A(n751), .Z(n588) );
  HS65_LL_AOI21X2 U583 ( .A(N210), .B(n732), .C(n731), .Z(n825) );
  HS65_LL_AOI21X2 U584 ( .A(N1138), .B(n943), .C(n971), .Z(n529) );
  HS65_LL_IVX18 U585 ( .A(N348), .Z(N1138) );
  HS65_LL_BFX35 U586 ( .A(N335), .Z(n819) );
  HS65_LL_NOR4ABX4 U587 ( .A(n987), .B(n986), .C(n985), .D(n984), .Z(n988) );
  HS65_LL_OR2X27 U588 ( .A(n1026), .B(n1025), .Z(N6926) );
  HS65_LL_OR2ABX18 U589 ( .A(n1059), .B(n1058), .Z(N7761) );
  HS65_LH_NAND2X2 U590 ( .A(n1138), .B(n1121), .Z(n1058) );
  HS65_LL_AOI12X2 U591 ( .A(n1136), .B(n1122), .C(n1057), .Z(n1059) );
  HS65_LH_IVX71 U592 ( .A(n485), .Z(N6716) );
  HS65_LH_IVX2 U593 ( .A(n710), .Z(n487) );
  HS65_LH_IVX71 U594 ( .A(n487), .Z(N4740) );
  HS65_LH_NOR2X2 U595 ( .A(n709), .B(n708), .Z(n710) );
  HS65_LH_IVX2 U596 ( .A(n704), .Z(n489) );
  HS65_LH_IVX71 U597 ( .A(n489), .Z(N4739) );
  HS65_LH_NOR2X2 U598 ( .A(n703), .B(n708), .Z(n704) );
  HS65_LH_IVX2 U599 ( .A(n702), .Z(n491) );
  HS65_LH_IVX71 U600 ( .A(n491), .Z(N4738) );
  HS65_LH_NOR2X2 U601 ( .A(n701), .B(n708), .Z(n702) );
  HS65_LH_IVX2 U602 ( .A(n706), .Z(n493) );
  HS65_LH_NOR2X2 U603 ( .A(n705), .B(n708), .Z(n706) );
  HS65_LL_NOR2AX19 U604 ( .A(N136), .B(N1066), .Z(N2054) );
  HS65_LH_IVX2 U605 ( .A(n695), .Z(n495) );
  HS65_LH_IVX2 U606 ( .A(n692), .Z(n497) );
  HS65_LH_OAI212X3 U607 ( .A(N588), .B(N86), .C(n707), .D(N87), .E(n1140), .Z(
        n692) );
  HS65_LH_IVX2 U608 ( .A(n513), .Z(n499) );
  HS65_LH_IVX71 U609 ( .A(n499), .Z(N6643) );
  HS65_LH_AND3X4 U610 ( .A(n997), .B(n674), .C(n503), .Z(n513) );
  HS65_LH_IVX2 U611 ( .A(n693), .Z(n501) );
  HS65_LH_IVX71 U612 ( .A(n501), .Z(N4278) );
  HS65_LH_OAI212X3 U613 ( .A(N588), .B(N88), .C(n707), .D(N34), .E(n1140), .Z(
        n693) );
  HS65_LH_MUXI41X2 U614 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(N265), .S1(N400), .Z(n864) );
  HS65_LHS_XNOR2X6 U615 ( .A(n867), .B(n866), .Z(n868) );
  HS65_LH_AOI12X3 U616 ( .A(n990), .B(n1020), .C(n820), .Z(n821) );
  HS65_LH_OR2X9 U617 ( .A(n943), .B(n536), .Z(n521) );
  HS65_LH_IVX9 U618 ( .A(n679), .Z(n682) );
  HS65_LHS_XNOR2X6 U619 ( .A(n610), .B(n609), .Z(n616) );
  HS65_LHS_XNOR2X6 U620 ( .A(n932), .B(n1017), .Z(n933) );
  HS65_LH_IVX9 U621 ( .A(n793), .Z(n681) );
  HS65_LH_IVX2 U622 ( .A(N54), .Z(n636) );
  HS65_LH_AOI22X11 U623 ( .A(n819), .B(n622), .C(n621), .D(n732), .Z(n803) );
  HS65_LH_NAND2X2 U624 ( .A(N53), .B(n1011), .Z(n884) );
  HS65_LH_MUXI21X15 U625 ( .D0(N361), .D1(N366), .S0(n943), .Z(n952) );
  HS65_LH_NAND2X14 U626 ( .A(n834), .B(n887), .Z(n841) );
  HS65_LH_NAND2X2 U627 ( .A(n1065), .B(n1068), .Z(n1066) );
  HS65_LH_XNOR2X9 U628 ( .A(n841), .B(n915), .Z(n900) );
  HS65_LH_AND2X4 U629 ( .A(n761), .B(n763), .Z(n1115) );
  HS65_LH_IVX2 U630 ( .A(n645), .Z(n643) );
  HS65_LH_IVX2 U631 ( .A(n831), .Z(n930) );
  HS65_LH_NAND2X2 U632 ( .A(N119), .B(n1011), .Z(n974) );
  HS65_LH_NAND2X14 U633 ( .A(n771), .B(n770), .Z(n1001) );
  HS65_LH_IVX2 U634 ( .A(N503), .Z(n585) );
  HS65_LH_NOR2X2 U635 ( .A(n990), .B(n1020), .Z(n991) );
  HS65_LH_NAND2X2 U636 ( .A(n1138), .B(n1075), .Z(n892) );
  HS65_LH_NAND2X14 U637 ( .A(n514), .B(n741), .Z(n1120) );
  HS65_LH_IVX2 U638 ( .A(N7473), .Z(n1123) );
  HS65_LH_IVX2 U639 ( .A(N210), .Z(n733) );
  HS65_LL_BFX9 U640 ( .A(n673), .Z(n503) );
  HS65_LL_IVX9 U641 ( .A(N341), .Z(n536) );
  HS65_LL_IVX18 U642 ( .A(n1161), .Z(n504) );
  HS65_LL_IVX27 U643 ( .A(n504), .Z(N8123) );
  HS65_LL_NAND2X7 U644 ( .A(n1056), .B(n1055), .Z(n1161) );
  HS65_LLS_XOR2X6 U645 ( .A(n956), .B(n591), .Z(n592) );
  HS65_LL_BFX53 U646 ( .A(N332), .Z(n943) );
  HS65_LLS_XNOR2X6 U647 ( .A(N273), .B(N411), .Z(n624) );
  HS65_LL_IVX9 U648 ( .A(n669), .Z(n670) );
  HS65_LL_NAND2X14 U649 ( .A(n522), .B(n1072), .Z(N8128) );
  HS65_LL_NAND2X7 U650 ( .A(n516), .B(n1038), .Z(n1085) );
  HS65_LH_IVX22 U651 ( .A(n1121), .Z(N7704) );
  HS65_LH_NAND2X7 U652 ( .A(n1128), .B(n1120), .Z(n742) );
  HS65_LH_NAND2X7 U653 ( .A(n1132), .B(n1122), .Z(n1091) );
  HS65_LH_NAND2X5 U654 ( .A(n1136), .B(n1114), .Z(n1061) );
  HS65_LH_NAND2X5 U655 ( .A(n1138), .B(n1060), .Z(n1062) );
  HS65_LH_IVX22 U656 ( .A(n1114), .Z(N7702) );
  HS65_LH_NAND2AX7 U657 ( .A(n779), .B(n778), .Z(n1060) );
  HS65_LL_NAND2X2 U658 ( .A(n847), .B(n844), .Z(n845) );
  HS65_LH_NOR2X6 U659 ( .A(n1037), .B(n1010), .Z(n1015) );
  HS65_LH_NOR2X6 U660 ( .A(n655), .B(n656), .Z(n657) );
  HS65_LH_NOR2X6 U661 ( .A(n904), .B(n993), .Z(n688) );
  HS65_LL_NOR2X5 U662 ( .A(n681), .B(n633), .Z(n656) );
  HS65_LH_NAND3X3 U663 ( .A(n715), .B(n753), .C(n580), .Z(n581) );
  HS65_LL_NAND2X4 U664 ( .A(n583), .B(n582), .Z(n584) );
  HS65_LH_NAND2X7 U665 ( .A(n1040), .B(n1035), .Z(n872) );
  HS65_LL_AO222X4 U666 ( .A(n697), .B(n1042), .C(n1011), .D(N129), .E(n1040), 
        .F(n985), .Z(n508) );
  HS65_LH_IVX7 U667 ( .A(n714), .Z(n580) );
  HS65_LL_OAI21X5 U668 ( .A(n785), .B(n511), .C(n515), .Z(n790) );
  HS65_LL_AOI12X4 U669 ( .A(n784), .B(n908), .C(n786), .Z(n633) );
  HS65_LH_OA12X9 U670 ( .A(n757), .B(n588), .C(n1117), .Z(n597) );
  HS65_LH_NAND2X7 U671 ( .A(n763), .B(n1117), .Z(n767) );
  HS65_LL_NAND2X5 U672 ( .A(n629), .B(n799), .Z(n908) );
  HS65_LH_NOR2AX3 U673 ( .A(N54), .B(n716), .Z(n717) );
  HS65_LH_NAND2X7 U674 ( .A(n777), .B(n776), .Z(n779) );
  HS65_LL_NOR2X3 U675 ( .A(n682), .B(n799), .Z(n687) );
  HS65_LH_AOI22X4 U676 ( .A(N173), .B(n1135), .C(N203), .D(n1134), .Z(n1063)
         );
  HS65_LL_OAI12X3 U677 ( .A(n506), .B(n982), .C(n974), .Z(n975) );
  HS65_LH_NAND2AX7 U678 ( .A(n801), .B(n630), .Z(n805) );
  HS65_LH_OAI21X6 U679 ( .A(n1037), .B(n755), .C(n672), .Z(n507) );
  HS65_LL_AOI12X4 U680 ( .A(n902), .B(n907), .C(n809), .Z(n799) );
  HS65_LH_NAND2X5 U681 ( .A(n679), .B(n655), .Z(n684) );
  HS65_LH_IVX2 U682 ( .A(n887), .Z(n838) );
  HS65_LH_IVX9 U683 ( .A(n638), .Z(n557) );
  HS65_LH_NAND2X4 U684 ( .A(n1040), .B(n1105), .Z(n776) );
  HS65_LH_IVX9 U685 ( .A(n576), .Z(n745) );
  HS65_LH_NOR2X5 U686 ( .A(n1008), .B(n506), .Z(n1016) );
  HS65_LH_NOR2X6 U687 ( .A(n1096), .B(n762), .Z(n769) );
  HS65_LH_NAND2X5 U688 ( .A(N112), .B(n1011), .Z(n780) );
  HS65_LH_OR2ABX27 U689 ( .A(n1140), .B(N140), .Z(N2590) );
  HS65_LH_OR2ABX27 U690 ( .A(n1140), .B(N83), .Z(N4279) );
  HS65_LH_IVX9 U691 ( .A(n928), .Z(n630) );
  HS65_LL_IVX4 U692 ( .A(n534), .Z(n949) );
  HS65_LL_NAND2X2 U693 ( .A(n585), .B(n950), .Z(n583) );
  HS65_LL_MUXI21X2 U694 ( .D0(N308), .D1(N315), .S0(n943), .Z(n947) );
  HS65_LH_IVX9 U695 ( .A(N595), .Z(n921) );
  HS65_LHS_XOR2X3 U696 ( .A(N341), .B(N351), .Z(n965) );
  HS65_LH_IVX22 U697 ( .A(N366), .Z(N1139) );
  HS65_LL_IVX18 U698 ( .A(N358), .Z(N1145) );
  HS65_LH_IVX7 U699 ( .A(N613), .Z(n725) );
  HS65_LL_NAND2X5 U700 ( .A(n1088), .B(n1087), .Z(n1089) );
  HS65_LL_NOR2AX3 U701 ( .A(n1069), .B(n1085), .Z(n1070) );
  HS65_LL_NAND2X5 U702 ( .A(n1128), .B(n1085), .Z(n1047) );
  HS65_LL_AOI12X4 U703 ( .A(N571), .B(n1085), .C(N574), .Z(n1088) );
  HS65_LH_NAND2X7 U704 ( .A(n1133), .B(n1120), .Z(n1032) );
  HS65_LL_OA12X9 U705 ( .A(n874), .B(n1041), .C(n523), .Z(n510) );
  HS65_LL_NAND2X14 U706 ( .A(n998), .B(n772), .Z(N7432) );
  HS65_LH_AOI12X6 U707 ( .A(n1132), .B(n1119), .C(n1031), .Z(n1033) );
  HS65_LL_OAI12X6 U708 ( .A(n1037), .B(n1005), .C(n512), .Z(n1121) );
  HS65_LH_NAND2X7 U709 ( .A(n913), .B(n912), .Z(n919) );
  HS65_LL_NAND2X4 U710 ( .A(n1042), .B(n899), .Z(n890) );
  HS65_LH_NOR3X2 U711 ( .A(n759), .B(n758), .C(n781), .Z(n773) );
  HS65_LH_IVX9 U712 ( .A(n1003), .Z(n1005) );
  HS65_LH_NAND2X7 U713 ( .A(n1042), .B(n774), .Z(n664) );
  HS65_LL_OAI21X3 U714 ( .A(n595), .B(n594), .C(n593), .Z(n596) );
  HS65_LH_NAND2X7 U715 ( .A(n1042), .B(n900), .Z(n778) );
  HS65_LH_NAND2X7 U716 ( .A(n1042), .B(n781), .Z(n782) );
  HS65_LLS_XNOR2X3 U717 ( .A(n740), .B(n739), .Z(n920) );
  HS65_LL_OAI12X3 U718 ( .A(n916), .B(n915), .C(n914), .Z(n917) );
  HS65_LL_NAND2X4 U719 ( .A(n570), .B(n567), .Z(n568) );
  HS65_LH_NAND2X5 U720 ( .A(n527), .B(n1021), .Z(n847) );
  HS65_LH_NAND2X7 U721 ( .A(n1042), .B(n910), .Z(n634) );
  HS65_LH_IVX9 U722 ( .A(N7467), .Z(n1137) );
  HS65_LH_NAND2X7 U723 ( .A(n544), .B(n661), .Z(n662) );
  HS65_LL_NAND2AX7 U724 ( .A(n688), .B(n1021), .Z(n915) );
  HS65_LL_NOR2X6 U725 ( .A(n996), .B(n719), .Z(n1116) );
  HS65_LL_OAI21X6 U726 ( .A(n950), .B(n585), .C(n584), .Z(n996) );
  HS65_LL_NOR2X3 U727 ( .A(n756), .B(n749), .Z(n719) );
  HS65_LH_NAND2X7 U728 ( .A(n769), .B(n768), .Z(n770) );
  HS65_LLS_XNOR2X3 U729 ( .A(n790), .B(n789), .Z(n796) );
  HS65_LH_IVX9 U730 ( .A(n767), .Z(n768) );
  HS65_LH_NAND2X4 U731 ( .A(n762), .B(n997), .Z(n722) );
  HS65_LH_NAND2X7 U732 ( .A(n718), .B(n717), .Z(n749) );
  HS65_LH_NAND2X7 U733 ( .A(n992), .B(n991), .Z(n1022) );
  HS65_LH_IVX9 U734 ( .A(n1009), .Z(n1010) );
  HS65_LH_IVX9 U735 ( .A(n798), .Z(n686) );
  HS65_LLS_XNOR2X3 U736 ( .A(n909), .B(n908), .Z(n1009) );
  HS65_LLS_XNOR2X3 U737 ( .A(n616), .B(n615), .Z(n1039) );
  HS65_LL_AOI21X2 U738 ( .A(n841), .B(n885), .C(n992), .Z(n822) );
  HS65_LH_IVX9 U739 ( .A(n555), .Z(n566) );
  HS65_LLS_XNOR2X3 U740 ( .A(n812), .B(n811), .Z(n813) );
  HS65_LL_NAND3X3 U741 ( .A(n684), .B(n683), .C(n517), .Z(n685) );
  HS65_LL_NAND2X4 U742 ( .A(n952), .B(n640), .Z(n714) );
  HS65_LH_NAND2X7 U743 ( .A(n793), .B(n784), .Z(n798) );
  HS65_LH_NOR2X6 U744 ( .A(n885), .B(n841), .Z(n992) );
  HS65_LH_NOR2X5 U745 ( .A(n805), .B(n681), .Z(n787) );
  HS65_LL_OAI21X2 U746 ( .A(n825), .B(n824), .C(n828), .Z(n826) );
  HS65_LH_AOI22X6 U747 ( .A(N167), .B(n1131), .C(N197), .D(n1130), .Z(n1073)
         );
  HS65_LH_IVX9 U748 ( .A(n834), .Z(n886) );
  HS65_LH_IVX9 U749 ( .A(n1106), .Z(n728) );
  HS65_LH_IVX9 U750 ( .A(n805), .Z(n786) );
  HS65_LL_OR2X4 U751 ( .A(n904), .B(n800), .Z(n629) );
  HS65_LH_IVX9 U752 ( .A(n800), .Z(n677) );
  HS65_LH_AOI22X6 U753 ( .A(N167), .B(n1135), .C(N197), .D(n1134), .Z(n879) );
  HS65_LL_NAND2X4 U754 ( .A(n546), .B(n557), .Z(n547) );
  HS65_LH_IVX9 U755 ( .A(n543), .Z(n544) );
  HS65_LH_IVX9 U756 ( .A(n763), .Z(n995) );
  HS65_LH_IVX9 U757 ( .A(n668), .Z(n666) );
  HS65_LH_IVX9 U758 ( .A(n994), .Z(n674) );
  HS65_LH_IVX9 U759 ( .A(n715), .Z(n663) );
  HS65_LH_NAND2AX7 U760 ( .A(n676), .B(n675), .Z(n834) );
  HS65_LH_IVX9 U761 ( .A(n1020), .Z(n918) );
  HS65_LH_NOR2X6 U762 ( .A(N374), .B(n808), .Z(n905) );
  HS65_LH_NAND2X7 U763 ( .A(n652), .B(n651), .Z(n791) );
  HS65_LHS_XNOR2X3 U764 ( .A(n934), .B(n933), .Z(n936) );
  HS65_LH_IVX9 U765 ( .A(n902), .Z(n903) );
  HS65_LL_NOR2X5 U766 ( .A(n535), .B(n949), .Z(n543) );
  HS65_LH_NAND2X7 U767 ( .A(n713), .B(n712), .Z(n724) );
  HS65_LH_IVX9 U768 ( .A(n1109), .Z(n1008) );
  HS65_LH_IVX9 U769 ( .A(n1011), .Z(n1012) );
  HS65_LH_NAND2X7 U770 ( .A(n636), .B(n952), .Z(n696) );
  HS65_LH_IVX4 U771 ( .A(n1125), .Z(n1054) );
  HS65_LL_NOR2X5 U772 ( .A(N534), .B(n953), .Z(n556) );
  HS65_LL_NAND2X5 U773 ( .A(N534), .B(n953), .Z(n552) );
  HS65_LH_NAND2X7 U774 ( .A(N116), .B(n1011), .Z(n876) );
  HS65_LH_NAND2X7 U775 ( .A(n732), .B(n650), .Z(n651) );
  HS65_LH_NAND2X7 U776 ( .A(n761), .B(n1096), .Z(n994) );
  HS65_LH_AND2ABX18 U777 ( .A(N580), .B(n667), .Z(n1138) );
  HS65_LL_NAND2X5 U778 ( .A(n734), .B(n934), .Z(n837) );
  HS65_LH_IVX9 U779 ( .A(n931), .Z(n675) );
  HS65_LH_NAND2X7 U780 ( .A(n676), .B(n931), .Z(n887) );
  HS65_LL_NAND2X4 U781 ( .A(N457), .B(n831), .Z(n828) );
  HS65_LH_IVX9 U782 ( .A(n680), .Z(n927) );
  HS65_LH_IVX9 U783 ( .A(N709), .Z(n708) );
  HS65_LH_IVX9 U784 ( .A(n999), .Z(n1098) );
  HS65_LH_NAND2X4 U785 ( .A(n1040), .B(n979), .Z(n712) );
  HS65_LH_NOR3X4 U786 ( .A(N1152), .B(N1155), .C(N2061), .Z(n969) );
  HS65_LH_NAND2X7 U787 ( .A(N2139), .B(N577), .Z(n667) );
  HS65_LH_NAND2X7 U788 ( .A(N2139), .B(N571), .Z(n644) );
  HS65_LH_IVX4 U789 ( .A(n1129), .Z(n895) );
  HS65_LH_AOI22X6 U790 ( .A(N103), .B(n1029), .C(N100), .D(n1124), .Z(n1048)
         );
  HS65_LH_IVX9 U791 ( .A(N583), .Z(n570) );
  HS65_LH_IVX9 U792 ( .A(N4), .Z(n904) );
  HS65_LH_IVX9 U793 ( .A(N389), .Z(n654) );
  HS65_LH_IVX9 U794 ( .A(N225), .Z(n735) );
  HS65_LH_IVX9 U795 ( .A(N468), .Z(n734) );
  HS65_LH_IVX9 U796 ( .A(N422), .Z(n676) );
  HS65_LH_IVX9 U797 ( .A(N596), .Z(n922) );
  HS65_LH_IVX9 U798 ( .A(N374), .Z(n626) );
  HS65_LH_IVX9 U799 ( .A(N446), .Z(n1018) );
  HS65_LH_IVX9 U800 ( .A(N479), .Z(n574) );
  HS65_LH_IVX9 U801 ( .A(N610), .Z(n1028) );
  HS65_LH_IVX9 U802 ( .A(N127), .Z(n1013) );
  HS65_LH_IVX9 U803 ( .A(N603), .Z(n1100) );
  HS65_LH_IVX9 U804 ( .A(N514), .Z(n535) );
  HS65_LH_IVX9 U805 ( .A(N490), .Z(n571) );
  HS65_LH_IVX9 U806 ( .A(N588), .Z(n707) );
  HS65_LLS_XNOR2X3 U807 ( .A(N288), .B(N374), .Z(n622) );
  HS65_LH_IVX9 U808 ( .A(N115), .Z(n1004) );
  HS65_LH_IVX9 U809 ( .A(N114), .Z(n729) );
  HS65_LHS_XOR2X6 U810 ( .A(N234), .B(N435), .Z(n650) );
  HS65_LL_NAND2X14 U811 ( .A(n1090), .B(n1089), .Z(N8127) );
  HS65_LL_NOR2X6 U812 ( .A(n1071), .B(n1070), .Z(n1072) );
  HS65_LL_AOI12X6 U813 ( .A(n1126), .B(n1086), .C(n1053), .Z(n1056) );
  HS65_LH_NAND2AX7 U814 ( .A(n1054), .B(n1085), .Z(n1055) );
  HS65_LL_AOI12X6 U815 ( .A(n1129), .B(n1086), .C(n1045), .Z(n1046) );
  HS65_LL_NAND2X7 U816 ( .A(n1044), .B(n1043), .Z(n1086) );
  HS65_LL_MUX21I1X6 U817 ( .D0(n1097), .D1(N7432), .S0(N599), .Z(n1102) );
  HS65_LH_IVX27 U818 ( .A(n510), .Z(N8075) );
  HS65_LL_NAND2X14 U819 ( .A(n1077), .B(n1076), .Z(N7755) );
  HS65_LL_NAND4ABX3 U820 ( .A(n774), .B(n878), .C(n773), .D(N7432), .Z(n775)
         );
  HS65_LL_NAND2X2 U821 ( .A(n1133), .B(n1121), .Z(n1092) );
  HS65_LH_NAND2X7 U822 ( .A(n1133), .B(n1075), .Z(n1076) );
  HS65_LH_NAND2X5 U823 ( .A(n1129), .B(n1119), .Z(n743) );
  HS65_LL_NAND2X5 U824 ( .A(n1042), .B(n1041), .Z(n1043) );
  HS65_LL_NAND2AX7 U825 ( .A(n1037), .B(n1036), .Z(n1038) );
  HS65_LH_NAND2X5 U826 ( .A(n1126), .B(n1079), .Z(n1080) );
  HS65_LL_NAND2AX7 U827 ( .A(n891), .B(n890), .Z(n1075) );
  HS65_LL_AOI12X6 U828 ( .A(n1042), .B(n878), .C(n877), .Z(n1049) );
  HS65_LH_NAND2AX7 U829 ( .A(n1037), .B(n920), .Z(n741) );
  HS65_LL_NAND2X4 U830 ( .A(n1042), .B(n758), .Z(n723) );
  HS65_LL_NOR3AX2 U831 ( .A(n901), .B(n900), .C(n899), .Z(n913) );
  HS65_LLS_XNOR2X6 U832 ( .A(n848), .B(n518), .Z(n849) );
  HS65_LL_AO222X4 U833 ( .A(n900), .B(n1042), .C(n1011), .D(N113), .E(n1040), 
        .F(n1105), .Z(n691) );
  HS65_LL_OAI211X3 U834 ( .A(n722), .B(n1116), .C(n721), .D(n720), .Z(n758) );
  HS65_LH_NAND2X5 U835 ( .A(n1125), .B(n1078), .Z(n1081) );
  HS65_LLS_XNOR2X3 U836 ( .A(n889), .B(n888), .Z(n899) );
  HS65_LL_AOI12X3 U837 ( .A(n887), .B(n915), .C(n886), .Z(n888) );
  HS65_LL_NAND2X4 U838 ( .A(n594), .B(n592), .Z(n593) );
  HS65_LH_NAND2X5 U839 ( .A(n1115), .B(n1116), .Z(n720) );
  HS65_LLS_XNOR2X3 U840 ( .A(n663), .B(n662), .Z(n774) );
  HS65_LL_NAND2X4 U841 ( .A(n640), .B(n639), .Z(n661) );
  HS65_LH_AOI21X6 U842 ( .A(n633), .B(n681), .C(n656), .Z(n910) );
  HS65_LL_AOI12X23 U843 ( .A(n1042), .B(n976), .C(n975), .Z(N7467) );
  HS65_LH_NOR2X5 U844 ( .A(n1022), .B(n1021), .Z(n1023) );
  HS65_LL_AOI21X4 U845 ( .A(n687), .B(n686), .C(n685), .Z(n1021) );
  HS65_LL_NAND2X4 U846 ( .A(n842), .B(n1019), .Z(n914) );
  HS65_LL_NOR2AX3 U847 ( .A(n715), .B(n714), .Z(n718) );
  HS65_LH_IVX9 U848 ( .A(n990), .Z(n740) );
  HS65_LH_NOR2X3 U849 ( .A(n990), .B(n1020), .Z(n820) );
  HS65_LH_NOR2X5 U850 ( .A(n1020), .B(n1019), .Z(n1024) );
  HS65_LL_NAND2AX7 U851 ( .A(n548), .B(n547), .Z(n582) );
  HS65_LH_IVX4 U852 ( .A(n558), .Z(n562) );
  HS65_LL_NAND2X5 U853 ( .A(n588), .B(n757), .Z(n1117) );
  HS65_LLS_XNOR2X3 U854 ( .A(n907), .B(n906), .Z(n926) );
  HS65_LH_NOR2X5 U855 ( .A(n787), .B(n655), .Z(n797) );
  HS65_LH_NOR2X3 U856 ( .A(n590), .B(n588), .Z(n589) );
  HS65_LLS_XNOR2X3 U857 ( .A(n940), .B(n939), .Z(n941) );
  HS65_LL_CBI4I1X3 U858 ( .A(n952), .B(n552), .C(n545), .D(n544), .Z(n548) );
  HS65_LH_OA22X9 U859 ( .A(n1012), .B(n729), .C(n506), .D(n728), .Z(n514) );
  HS65_LL_AOI13X4 U860 ( .A(n886), .B(n827), .C(n837), .D(n826), .Z(n1019) );
  HS65_LH_NOR2X3 U861 ( .A(n557), .B(n952), .Z(n558) );
  HS65_LH_OAI211X3 U862 ( .A(n807), .B(n806), .C(n805), .D(n804), .Z(n812) );
  HS65_LLS_XNOR2X3 U863 ( .A(n936), .B(n935), .Z(n940) );
  HS65_LL_NOR2AX6 U864 ( .A(n546), .B(n543), .Z(n640) );
  HS65_LL_NAND2X4 U865 ( .A(n542), .B(n546), .Z(n545) );
  HS65_LH_OA12X9 U866 ( .A(n907), .B(n803), .C(n800), .Z(n792) );
  HS65_LL_NOR2X5 U867 ( .A(n747), .B(n745), .Z(n757) );
  HS65_LH_AOI22X4 U868 ( .A(N161), .B(n1131), .C(N191), .D(n1130), .Z(n1093)
         );
  HS65_LL_IVX7 U869 ( .A(n909), .Z(n784) );
  HS65_LL_NAND2AX7 U870 ( .A(n637), .B(n561), .Z(n756) );
  HS65_LL_NAND2X7 U871 ( .A(n803), .B(n907), .Z(n800) );
  HS65_LLS_XNOR2X3 U872 ( .A(n865), .B(n864), .Z(n866) );
  HS65_LH_OA22X9 U873 ( .A(n1103), .B(n506), .C(n1004), .D(n1012), .Z(n512) );
  HS65_LL_NAND2X7 U874 ( .A(n541), .B(n638), .Z(n716) );
  HS65_LH_AOI22X4 U875 ( .A(n1011), .B(N126), .C(n1040), .D(n1110), .Z(n925)
         );
  HS65_LL_IVX4 U876 ( .A(n556), .Z(n561) );
  HS65_LL_IVX7 U877 ( .A(n552), .Z(n637) );
  HS65_LL_AOI12X6 U878 ( .A(n747), .B(n588), .C(n586), .Z(n763) );
  HS65_LH_NOR2X5 U879 ( .A(n1013), .B(n1012), .Z(n1014) );
  HS65_LH_NAND2X5 U880 ( .A(N52), .B(n1011), .Z(n660) );
  HS65_LLS_XNOR2X3 U881 ( .A(n859), .B(n1103), .Z(n867) );
  HS65_LL_NAND2X4 U882 ( .A(n571), .B(n520), .Z(n576) );
  HS65_LH_NAND2X4 U883 ( .A(N113), .B(n1011), .Z(n777) );
  HS65_LH_IVX9 U884 ( .A(n761), .Z(n762) );
  HS65_LH_IVX7 U885 ( .A(n1096), .Z(n760) );
  HS65_LH_AOI22X4 U886 ( .A(N131), .B(n1011), .C(n1040), .D(n977), .Z(n672) );
  HS65_LH_AOI22X4 U887 ( .A(N103), .B(n711), .C(N100), .D(n1127), .Z(n894) );
  HS65_LH_AOI22X4 U888 ( .A(n1011), .B(N123), .C(n1040), .D(n1098), .Z(n1000)
         );
  HS65_LHS_XOR2X3 U889 ( .A(N132), .B(n1096), .Z(n1097) );
  HS65_LHS_XNOR2X6 U890 ( .A(N503), .B(n950), .Z(n715) );
  HS65_LH_NOR2AX13 U891 ( .A(N580), .B(n667), .Z(n1135) );
  HS65_LH_NAND3X5 U892 ( .A(N468), .B(n737), .C(n736), .Z(n824) );
  HS65_LL_NAND2AX4 U893 ( .A(n680), .B(n678), .Z(n679) );
  HS65_LH_NOR2X6 U894 ( .A(n654), .B(n653), .Z(n655) );
  HS65_LH_NAND2X5 U895 ( .A(N435), .B(n680), .Z(n683) );
  HS65_LL_AOI22X6 U896 ( .A(n819), .B(n625), .C(n732), .D(n624), .Z(n907) );
  HS65_LH_IVX4 U897 ( .A(n932), .Z(n808) );
  HS65_LH_NOR2X5 U898 ( .A(n1018), .B(n1017), .Z(n1026) );
  HS65_LL_MUXI21X2 U899 ( .D0(N816), .D1(N299), .S0(n943), .Z(n1096) );
  HS65_LLS_XNOR2X3 U900 ( .A(N272), .B(n801), .Z(n620) );
  HS65_LL_MUXI21X2 U901 ( .D0(N302), .D1(N307), .S0(n943), .Z(n761) );
  HS65_LL_MUXI21X5 U902 ( .D0(N324), .D1(N331), .S0(n943), .Z(n950) );
  HS65_LH_NAND2X5 U903 ( .A(n819), .B(n649), .Z(n652) );
  HS65_LH_NOR2X3 U904 ( .A(n819), .B(N273), .Z(n627) );
  HS65_LL_NAND2AX4 U905 ( .A(N338), .B(n943), .Z(n534) );
  HS65_LL_MUXI21X2 U906 ( .D0(N226), .D1(N233), .S0(n819), .Z(n931) );
  HS65_LH_NAND2X5 U907 ( .A(N468), .B(n881), .Z(n882) );
  HS65_LH_NAND2X5 U908 ( .A(n819), .B(N217), .Z(n730) );
  HS65_LH_NOR2AX6 U909 ( .A(N616), .B(N613), .Z(n1127) );
  HS65_LH_NAND2AX29 U910 ( .A(N591), .B(N27), .Z(N2060) );
  HS65_LH_IVX9 U911 ( .A(N351), .Z(n611) );
  HS65_LH_IVX7 U912 ( .A(N411), .Z(n623) );
  HS65_LHS_XOR2X6 U913 ( .A(N241), .B(N435), .Z(n649) );
  HS65_LH_IVX7 U914 ( .A(N251), .Z(n858) );
  HS65_LH_IVX7 U915 ( .A(N435), .Z(n678) );
  HS65_LLS_XNOR2X3 U916 ( .A(N264), .B(N389), .Z(n632) );
  HS65_LH_IVX7 U917 ( .A(N566), .Z(n823) );
  HS65_LH_IVX27 U918 ( .A(n775), .Z(N7504) );
  HS65_LL_AOI12X23 U919 ( .A(N603), .B(n1102), .C(n1101), .Z(N7626) );
  HS65_LH_OR2X27 U920 ( .A(n1052), .B(n1051), .Z(N7738) );
  HS65_LL_BFX18 U921 ( .A(n875), .Z(N8076) );
  HS65_LL_IVX7 U922 ( .A(n646), .Z(n647) );
  HS65_LL_NAND2AX14 U923 ( .A(n893), .B(n892), .Z(N7759) );
  HS65_LL_OR3ABCX18 U924 ( .A(n1093), .B(n1092), .C(n1091), .Z(N7757) );
  HS65_LL_NAND2AX14 U925 ( .A(n897), .B(n896), .Z(N7741) );
  HS65_LH_IVX22 U926 ( .A(n1075), .Z(N7706) );
  HS65_LL_MX41X14 U927 ( .D0(n1119), .S0(n1126), .D1(n1120), .S1(n1125), .D2(
        n1029), .S2(N49), .D3(n1124), .S3(N46), .Z(N7737) );
  HS65_LL_MX41X14 U928 ( .D0(n1122), .S0(n1126), .D1(n1121), .S1(n1125), .D2(
        n1029), .S2(N106), .D3(n1124), .S3(N109), .Z(N7736) );
  HS65_LL_MX41X4 U929 ( .D0(n1064), .S0(n1138), .D1(n1030), .S1(n1136), .D2(
        n1135), .S2(N146), .D3(n1134), .S3(N149), .Z(n669) );
  HS65_LH_IVX22 U930 ( .A(n1120), .Z(N7705) );
  HS65_LL_OA12X9 U931 ( .A(n1074), .B(N7701), .C(n1073), .Z(n1077) );
  HS65_LL_MX41X14 U932 ( .D0(n1030), .S0(n1126), .D1(n1064), .S1(n1125), .D2(
        n1029), .S2(N20), .D3(n1124), .S3(N76), .Z(N7516) );
  HS65_LH_IVX22 U933 ( .A(n1119), .Z(N7700) );
  HS65_LL_OR3ABCX18 U934 ( .A(n1063), .B(n1062), .C(n1061), .Z(N7758) );
  HS65_LL_AND2X4 U935 ( .A(n1125), .B(n1075), .Z(n1051) );
  HS65_LH_MX41X7 U936 ( .D0(n1064), .S0(n1133), .D1(n1030), .S1(n1132), .D2(
        n1131), .S2(N146), .D3(n1130), .S3(N149), .Z(n646) );
  HS65_LH_IVX22 U937 ( .A(n1079), .Z(N7465) );
  HS65_LL_IVX7 U938 ( .A(N7466), .Z(n1030) );
  HS65_LL_NAND2AX7 U939 ( .A(n724), .B(n723), .Z(n1119) );
  HS65_LLS_XNOR2X6 U940 ( .A(n599), .B(n598), .Z(n1041) );
  HS65_LL_OAI12X3 U941 ( .A(n1050), .B(n1049), .C(n1048), .Z(n1052) );
  HS65_LH_IVX22 U942 ( .A(n691), .Z(N7707) );
  HS65_LL_OAI12X2 U943 ( .A(n880), .B(n1049), .C(n879), .Z(n893) );
  HS65_LH_IVX9 U944 ( .A(n1001), .Z(n772) );
  HS65_LLS_XNOR2X6 U945 ( .A(n850), .B(n849), .Z(n1036) );
  HS65_LLS_XNOR2X6 U946 ( .A(n597), .B(n596), .Z(n598) );
  HS65_LL_OA12X4 U947 ( .A(n1116), .B(n766), .C(n765), .Z(n771) );
  HS65_LL_OA12X4 U948 ( .A(n847), .B(n846), .C(n845), .Z(n518) );
  HS65_LLS_XNOR2X6 U949 ( .A(n751), .B(n526), .Z(n878) );
  HS65_LLS_XNOR2X3 U950 ( .A(n918), .B(n917), .Z(n1003) );
  HS65_LL_OAI12X6 U951 ( .A(n1037), .B(n754), .C(n641), .Z(n642) );
  HS65_LL_OAI21X2 U952 ( .A(n750), .B(n749), .C(n748), .Z(n526) );
  HS65_LH_NAND2AX7 U953 ( .A(n635), .B(n634), .Z(n1064) );
  HS65_LL_MUX21I1X6 U954 ( .D0(n818), .D1(n817), .S0(N566), .Z(n850) );
  HS65_LH_OR2X9 U955 ( .A(n1024), .B(n1023), .Z(n1025) );
  HS65_LLS_XNOR2X3 U956 ( .A(n791), .B(n657), .Z(n898) );
  HS65_LLS_XNOR2X3 U957 ( .A(n566), .B(n565), .Z(n567) );
  HS65_LL_OR2X4 U958 ( .A(n1015), .B(n1014), .Z(n519) );
  HS65_LHS_XNOR2X6 U959 ( .A(n551), .B(n550), .Z(n569) );
  HS65_LLS_XNOR2X3 U960 ( .A(n843), .B(n914), .Z(n844) );
  HS65_LLS_XNOR2X3 U961 ( .A(n579), .B(n578), .Z(n595) );
  HS65_LL_MX41X14 U962 ( .D0(n508), .S0(n1126), .D1(n1123), .S1(n1125), .D2(
        n1029), .S2(N70), .D3(n1124), .S3(N67), .Z(N7518) );
  HS65_LH_OR2X4 U963 ( .A(n823), .B(n993), .Z(n527) );
  HS65_LH_AOI31X3 U964 ( .A(n640), .B(n746), .C(n638), .D(n563), .Z(n550) );
  HS65_LLS_XNOR2X3 U965 ( .A(n564), .B(n563), .Z(n565) );
  HS65_LLS_XNOR2X3 U966 ( .A(n816), .B(n815), .Z(n817) );
  HS65_LH_IVX4 U967 ( .A(n1019), .Z(n916) );
  HS65_LH_OA22X9 U968 ( .A(n618), .B(n617), .C(n506), .D(n1039), .Z(n523) );
  HS65_LH_OA12X9 U969 ( .A(n506), .B(n1035), .C(n1034), .Z(n516) );
  HS65_LH_IVX27 U970 ( .A(n700), .Z(N7365) );
  HS65_LH_AOI22X4 U971 ( .A(N94), .B(N625), .C(n1040), .D(n1039), .Z(n1044) );
  HS65_LL_OAI12X3 U972 ( .A(n716), .B(n752), .C(n638), .Z(n639) );
  HS65_LLS_XNOR2X6 U973 ( .A(n753), .B(n752), .Z(n976) );
  HS65_LL_NAND3X5 U974 ( .A(n791), .B(n677), .C(n686), .Z(n993) );
  HS65_LLS_XNOR2X6 U975 ( .A(n814), .B(n813), .Z(n816) );
  HS65_LLS_XNOR2X3 U976 ( .A(n871), .B(n870), .Z(n1035) );
  HS65_LH_OR3X4 U977 ( .A(n990), .B(n841), .C(n885), .Z(n842) );
  HS65_LL_OA112X4 U978 ( .A(n562), .B(n561), .C(n560), .D(n559), .Z(n564) );
  HS65_LHS_XOR2X6 U979 ( .A(n696), .B(n746), .Z(n697) );
  HS65_LH_IVX9 U980 ( .A(n829), .Z(n738) );
  HS65_LLS_XNOR2X3 U981 ( .A(n532), .B(n531), .Z(n551) );
  HS65_LLS_XOR2X3 U982 ( .A(n797), .B(n799), .Z(n788) );
  HS65_LL_AOI12X4 U983 ( .A(n696), .B(n746), .C(n637), .Z(n752) );
  HS65_LH_IVX9 U984 ( .A(n756), .Z(n746) );
  HS65_LHS_XNOR2X3 U985 ( .A(n715), .B(n554), .Z(n555) );
  HS65_LH_NAND2X5 U986 ( .A(n1042), .B(n998), .Z(n1002) );
  HS65_LLS_XNOR2X3 U987 ( .A(n869), .B(n868), .Z(n870) );
  HS65_LH_IVX4 U988 ( .A(n1132), .Z(n1074) );
  HS65_LH_IVX4 U989 ( .A(n1136), .Z(n880) );
  HS65_LH_IVX9 U990 ( .A(n640), .Z(n549) );
  HS65_LH_AOI12X6 U991 ( .A(n837), .B(n886), .C(n839), .Z(n829) );
  HS65_LLS_XNOR2X3 U992 ( .A(n955), .B(n954), .Z(n957) );
  HS65_LH_IVX27 U993 ( .A(n507), .Z(N7015) );
  HS65_LH_NAND4ABX3 U994 ( .A(n1106), .B(n1105), .C(n1104), .D(n1103), .Z(
        n1112) );
  HS65_LL_CB4I6X4 U995 ( .A(n909), .B(n806), .C(n805), .D(n902), .Z(n515) );
  HS65_LLS_XNOR2X3 U996 ( .A(n854), .B(n853), .Z(n871) );
  HS65_LH_NAND2X4 U997 ( .A(n763), .B(n769), .Z(n764) );
  HS65_LH_OAI12X3 U998 ( .A(n905), .B(n904), .C(n903), .Z(n906) );
  HS65_LLS_XNOR2X3 U999 ( .A(n909), .B(n791), .Z(n795) );
  HS65_LL_MUXI21X2 U1000 ( .D0(n840), .D1(n839), .S0(n838), .Z(n843) );
  HS65_LH_IVX9 U1001 ( .A(n716), .Z(n753) );
  HS65_LH_MUXI21X2 U1002 ( .D0(n586), .D1(n577), .S0(n576), .Z(n525) );
  HS65_LH_OR3X4 U1003 ( .A(n682), .B(n681), .C(n805), .Z(n517) );
  HS65_LL_NAND2X4 U1004 ( .A(n762), .B(n587), .Z(n590) );
  HS65_LH_AOI21X2 U1005 ( .A(n952), .B(n556), .C(n553), .Z(n554) );
  HS65_LLS_XNOR2X3 U1006 ( .A(n606), .B(n605), .Z(n610) );
  HS65_LH_AO22X9 U1007 ( .A(N164), .B(n1131), .C(N194), .D(n1130), .Z(n1031)
         );
  HS65_LH_AO22X9 U1008 ( .A(N161), .B(n1135), .C(N191), .D(n1134), .Z(n1057)
         );
  HS65_LL_OAI22X4 U1009 ( .A(n620), .B(n732), .C(n619), .D(n937), .Z(n909) );
  HS65_LH_OAI12X3 U1010 ( .A(n506), .B(n986), .C(n660), .Z(n665) );
  HS65_LH_OAI211X1 U1011 ( .A(n808), .B(n803), .C(n907), .D(n802), .Z(n804) );
  HS65_LH_AO22X9 U1012 ( .A(N631), .B(N135), .C(n1100), .D(n1099), .Z(n1101)
         );
  HS65_LL_NAND2X5 U1013 ( .A(n837), .B(n824), .Z(n885) );
  HS65_LLS_XNOR2X3 U1014 ( .A(n603), .B(n602), .Z(n606) );
  HS65_LHS_XOR2X6 U1015 ( .A(n928), .B(n927), .Z(n929) );
  HS65_LHS_XNOR2X6 U1016 ( .A(n959), .B(n958), .Z(n964) );
  HS65_LH_IVX4 U1017 ( .A(n586), .Z(n587) );
  HS65_LL_AND2X4 U1018 ( .A(n541), .B(n540), .Z(n542) );
  HS65_LH_NAND3X3 U1019 ( .A(n983), .B(n982), .C(n981), .Z(n984) );
  HS65_LH_OAI12X3 U1020 ( .A(n506), .B(n1104), .C(n884), .Z(n891) );
  HS65_LH_OAI12X3 U1021 ( .A(n506), .B(n987), .C(n876), .Z(n877) );
  HS65_LH_MUX21I1X6 U1022 ( .D0(n727), .D1(n726), .S0(n832), .Z(n1106) );
  HS65_LHS_XNOR2X6 U1023 ( .A(N4), .B(n803), .Z(n911) );
  HS65_LH_OAI12X3 U1024 ( .A(n506), .B(n983), .C(n780), .Z(n783) );
  HS65_LH_NOR2X3 U1025 ( .A(n952), .B(n552), .Z(n553) );
  HS65_LL_AOI22X4 U1026 ( .A(n819), .B(n632), .C(n631), .D(n732), .Z(n793) );
  HS65_LH_AOI22X3 U1027 ( .A(N43), .B(n1124), .C(N37), .D(n1029), .Z(n1082) );
  HS65_LH_AOI22X4 U1028 ( .A(n1011), .B(N130), .C(n1040), .D(n978), .Z(n641)
         );
  HS65_LL_NOR2X5 U1029 ( .A(n574), .B(n947), .Z(n586) );
  HS65_LHS_XNOR2X6 U1030 ( .A(N54), .B(n952), .Z(n755) );
  HS65_LH_MUXI21X2 U1031 ( .D0(N251), .D1(N248), .S0(N210), .Z(n851) );
  HS65_LH_IVX9 U1032 ( .A(n732), .Z(n937) );
  HS65_LL_NOR2X5 U1033 ( .A(n571), .B(n520), .Z(n747) );
  HS65_LH_AO22X9 U1034 ( .A(N64), .B(n711), .C(N14), .D(n1127), .Z(n1045) );
  HS65_LH_NOR2AX13 U1035 ( .A(N574), .B(n644), .Z(n1131) );
  HS65_LL_NAND2X5 U1036 ( .A(n521), .B(n537), .Z(n541) );
  HS65_LLS_XNOR2X3 U1037 ( .A(n856), .B(n855), .Z(n869) );
  HS65_LL_NOR2X5 U1038 ( .A(n626), .B(n932), .Z(n902) );
  HS65_LH_OAI211X4 U1039 ( .A(n943), .B(n611), .C(n539), .D(n538), .Z(n540) );
  HS65_LH_NAND2X4 U1040 ( .A(N121), .B(n1011), .Z(n713) );
  HS65_LL_NAND2X5 U1041 ( .A(n509), .B(n535), .Z(n546) );
  HS65_LHS_XNOR2X6 U1042 ( .A(N210), .B(N218), .Z(n958) );
  HS65_LLS_XNOR2X3 U1043 ( .A(n861), .B(n860), .Z(n865) );
  HS65_LH_AO22X9 U1044 ( .A(N64), .B(n1029), .C(N14), .D(n1124), .Z(n1053) );
  HS65_LH_AOI22X3 U1045 ( .A(N49), .B(n711), .C(N46), .D(n1127), .Z(n744) );
  HS65_LL_NAND2X5 U1046 ( .A(n529), .B(n528), .Z(n638) );
  HS65_LL_AOI211X3 U1047 ( .A(n819), .B(n628), .C(n623), .D(n627), .Z(n809) );
  HS65_LHS_XNOR2X6 U1048 ( .A(n761), .B(n1096), .Z(n956) );
  HS65_LL_OR2X4 U1049 ( .A(n819), .B(N218), .Z(n736) );
  HS65_LH_AOI212X4 U1050 ( .A(N23), .B(N588), .C(N79), .D(n707), .E(N2623), 
        .Z(n703) );
  HS65_LL_MUXI21X2 U1051 ( .D0(N281), .D1(N288), .S0(n819), .Z(n932) );
  HS65_LH_MUX21I1X6 U1052 ( .D0(n659), .D1(n658), .S0(N503), .Z(n986) );
  HS65_LL_MUXI21X5 U1053 ( .D0(N265), .D1(N272), .S0(n819), .Z(n928) );
  HS65_LH_IVX4 U1054 ( .A(n1126), .Z(n1050) );
  HS65_LLS_XNOR2X3 U1055 ( .A(N265), .B(n801), .Z(n619) );
  HS65_LH_AOI212X4 U1056 ( .A(N25), .B(N588), .C(N24), .D(n707), .E(N2623), 
        .Z(n705) );
  HS65_LH_AOI212X4 U1057 ( .A(N81), .B(N588), .C(N26), .D(n707), .E(N2623), 
        .Z(n701) );
  HS65_LH_AOI212X4 U1058 ( .A(N80), .B(N588), .C(N82), .D(n707), .E(N2623), 
        .Z(n709) );
  HS65_LH_IVX18 U1059 ( .A(n819), .Z(n732) );
  HS65_LH_NAND2X5 U1060 ( .A(n943), .B(N358), .Z(n538) );
  HS65_LL_MUX41X9 U1061 ( .D0(n863), .D1(N251), .D2(n862), .D3(N248), .S0(N446), .S1(N206), .Z(n1103) );
  HS65_LH_IVX22 U1062 ( .A(N2527), .Z(N3613) );
  HS65_LH_MUX21I1X6 U1063 ( .D0(n733), .D1(N217), .S0(n819), .Z(n831) );
  HS65_LHS_XNOR2X6 U1064 ( .A(N292), .B(N264), .Z(n938) );
  HS65_LH_NOR2X2 U1065 ( .A(N120), .B(N619), .Z(n617) );
  HS65_LHS_XNOR2X6 U1066 ( .A(N372), .B(N323), .Z(n944) );
  HS65_LH_MUXI21X2 U1067 ( .D0(N597), .D1(N598), .S0(N226), .Z(n689) );
  HS65_LH_IVX4 U1068 ( .A(N280), .Z(n628) );
  HS65_LH_IVX7 U1069 ( .A(N534), .Z(n539) );
  HS65_LH_IVX22 U1070 ( .A(N552), .Z(N1153) );
  HS65_LH_IVX22 U1071 ( .A(N562), .Z(N1154) );
  HS65_LL_BFX62 U1072 ( .A(N1), .Z(N2309) );
  HS65_LHS_XNOR2X6 U1073 ( .A(N265), .B(N281), .Z(n959) );
  HS65_LHS_XNOR2X6 U1074 ( .A(N273), .B(N234), .Z(n962) );
  HS65_LHS_XNOR2X6 U1075 ( .A(N289), .B(N257), .Z(n961) );
  HS65_LLS_XNOR2X3 U1076 ( .A(N281), .B(N374), .Z(n621) );
  HS65_LH_IVX4 U1077 ( .A(N577), .Z(n1068) );
  HS65_LHS_XNOR2X6 U1078 ( .A(N226), .B(N206), .Z(n960) );
  HS65_LL_NAND2X14 U1079 ( .A(N386), .B(N556), .Z(N2061) );
  HS65_LL_NAND2X14 U1080 ( .A(N27), .B(N31), .Z(N2623) );
  HS65_LHS_XNOR2X6 U1081 ( .A(N257), .B(N389), .Z(n631) );
  HS65_LL_MX41X14 U1082 ( .D0(n1060), .S0(n1133), .D1(n1114), .S1(n1132), .D2(
        n1131), .S2(N173), .D3(n1130), .S3(N203), .Z(N7754) );
  HS65_LL_MUX21X4 U1083 ( .D0(n573), .D1(n572), .S0(n943), .Z(n751) );
  HS65_LL_MUXI21X5 U1084 ( .D0(n611), .D1(N1145), .S0(n943), .Z(n953) );
  HS65_LL_MUXI21X2 U1085 ( .D0(N316), .D1(N323), .S0(n943), .Z(n520) );
  HS65_LL_NAND2X14 U1086 ( .A(n1033), .B(n1032), .Z(N7756) );
  HS65_LL_MUX21X4 U1087 ( .D0(n836), .D1(n835), .S0(n834), .Z(n846) );
  HS65_LL_MX41X14 U1088 ( .D0(n1078), .S0(n1138), .D1(n1079), .S1(n1136), .D2(
        n1135), .S2(N170), .D3(n1134), .S3(N200), .Z(N7604) );
  HS65_LL_OR3ABCX18 U1089 ( .A(n1082), .B(n1081), .C(n1080), .Z(N7515) );
  HS65_LL_MX41X14 U1090 ( .D0(n1120), .S0(n1138), .D1(n1119), .S1(n1136), .D2(
        n1135), .S2(N164), .D3(n1134), .S3(N194), .Z(N7760) );
  HS65_LL_OA12X18 U1091 ( .A(n1037), .B(n926), .C(n925), .Z(N7473) );
  HS65_LL_MUXI21X2 U1092 ( .D0(n1019), .D1(n830), .S0(n829), .Z(n836) );
  HS65_LL_MX41X14 U1093 ( .D0(n1114), .S0(n1126), .D1(n1060), .S1(n1125), .D2(
        n1029), .S2(N40), .D3(n1124), .S3(N91), .Z(N7739) );
  HS65_LHS_XNOR2X6 U1094 ( .A(n795), .B(n794), .Z(n815) );
  HS65_LH_NAND2X2 U1095 ( .A(N97), .B(N625), .Z(n1034) );
  HS65_LH_NOR2X2 U1096 ( .A(N523), .B(n948), .Z(n530) );
  HS65_LHS_XNOR2X6 U1097 ( .A(n1018), .B(n1017), .Z(n1020) );
  HS65_LH_IVX2 U1098 ( .A(N580), .Z(n1065) );
  HS65_LH_NOR2X2 U1099 ( .A(N580), .B(n1068), .Z(n1069) );
  HS65_LL_NAND2AX7 U1100 ( .A(N571), .B(n1086), .Z(n1087) );
  HS65_LH_NAND2X2 U1101 ( .A(n576), .B(n746), .Z(n750) );
  HS65_LH_AOI12X2 U1102 ( .A(n576), .B(n996), .C(n747), .Z(n748) );
  HS65_LHS_XNOR2X3 U1103 ( .A(N369), .B(N316), .Z(n945) );
  HS65_LH_AO22X9 U1104 ( .A(N128), .B(n1011), .C(n1040), .D(n1107), .Z(n635)
         );
  HS65_LH_NOR2AX6 U1105 ( .A(N607), .B(N610), .Z(n1124) );
  HS65_LH_MUXI31X2 U1106 ( .D0(N596), .D1(N595), .D2(n698), .S0(N281), .S1(
        N374), .Z(n1113) );
  HS65_LH_IVX2 U1107 ( .A(n977), .Z(n980) );
  HS65_LH_MUXI41X2 U1108 ( .D0(N596), .D1(n1007), .D2(N595), .D3(n1006), .S0(
        N534), .S1(N351), .Z(n985) );
  HS65_LH_NAND2X2 U1109 ( .A(n801), .B(n928), .Z(n802) );
  HS65_LH_MUXI41X4 U1110 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(
        N234), .S1(N435), .Z(n860) );
  HS65_LH_MUXI41X4 U1111 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(
        N281), .S1(N374), .Z(n861) );
  HS65_LH_IVX2 U1112 ( .A(n809), .Z(n806) );
  HS65_LH_IVX2 U1113 ( .A(n802), .Z(n807) );
  HS65_LH_NOR2X2 U1114 ( .A(N411), .B(n935), .Z(n810) );
  HS65_LH_NAND2X2 U1115 ( .A(n832), .B(n930), .Z(n833) );
  HS65_LH_IVX2 U1116 ( .A(n828), .Z(n830) );
  HS65_LH_IVX2 U1117 ( .A(n837), .Z(n840) );
  HS65_LH_NAND2X2 U1118 ( .A(n902), .B(n805), .Z(n785) );
  HS65_LH_AOI22X1 U1119 ( .A(n557), .B(n952), .C(n716), .D(n558), .Z(n560) );
  HS65_LH_MUXI21X2 U1120 ( .D0(n590), .D1(n589), .S0(n747), .Z(n591) );
  HS65_LH_AOI12X2 U1121 ( .A(N583), .B(n503), .C(n996), .Z(n594) );
  HS65_LHS_XNOR2X3 U1122 ( .A(n1096), .B(n525), .Z(n579) );
  HS65_LH_NOR2X2 U1123 ( .A(N479), .B(n575), .Z(n577) );
  HS65_LH_MUXI41X2 U1124 ( .D0(N254), .D1(n858), .D2(N242), .D3(n857), .S0(
        N468), .S1(N218), .Z(n855) );
  HS65_LH_MUXI41X2 U1125 ( .D0(N254), .D1(n858), .D2(N242), .D3(n857), .S0(
        N422), .S1(N226), .Z(n856) );
  HS65_LH_NAND2X2 U1126 ( .A(n761), .B(n767), .Z(n578) );
  HS65_LHS_XNOR2X3 U1127 ( .A(n952), .B(n756), .Z(n532) );
  HS65_LHS_XNOR2X3 U1128 ( .A(n977), .B(n604), .Z(n605) );
  HS65_LH_MUXI21X2 U1129 ( .D0(N218), .D1(N225), .S0(n819), .Z(n934) );
  HS65_LHS_XNOR2X6 U1130 ( .A(N280), .B(N411), .Z(n625) );
  HS65_LH_NAND2X2 U1131 ( .A(n1096), .B(n997), .Z(n766) );
  HS65_LH_NAND2AX4 U1132 ( .A(n764), .B(n1116), .Z(n765) );
  HS65_LH_IVX9 U1133 ( .A(N242), .Z(n862) );
  HS65_LH_IVX2 U1134 ( .A(n898), .Z(n901) );
  HS65_LHS_XNOR2X6 U1135 ( .A(n968), .B(n967), .Z(n1094) );
  HS65_LH_AO12X4 U1136 ( .A(N580), .B(n1067), .C(n1083), .Z(n1071) );
  HS65_LH_AOI21X2 U1137 ( .A(N574), .B(n1084), .C(n1083), .Z(n1090) );
  HS65_LL_OAI112X1 U1138 ( .A(n874), .B(n1036), .C(n873), .D(n872), .Z(n875)
         );
  HS65_LH_BFX27 U1139 ( .A(n1049), .Z(N7701) );
  HS65_LH_XOR2X27 U1140 ( .A(N132), .B(n1118), .Z(N7698) );
  HS65_LH_IVX22 U1141 ( .A(n670), .Z(N7607) );
  HS65_LH_IVX27 U1142 ( .A(n647), .Z(N7603) );
  HS65_LH_XNOR2X27 U1143 ( .A(n957), .B(n956), .Z(N7474) );
  HS65_LH_IVX27 U1144 ( .A(n1064), .Z(N7471) );
  HS65_LH_IVX22 U1145 ( .A(n1078), .Z(N7470) );
  HS65_LH_IVX27 U1146 ( .A(n642), .Z(N7466) );
  HS65_LH_IVX27 U1147 ( .A(n508), .Z(N7363) );
  HS65_LH_XNOR2X27 U1148 ( .A(n964), .B(n963), .Z(N6877) );
  HS65_LH_AND3ABCX27 U1149 ( .A(n1113), .B(n1112), .C(n1111), .Z(N5388) );
  HS65_LH_BFX27 U1150 ( .A(N137), .Z(N2139) );
  HS65_LH_AND2X27 U1151 ( .A(N2309), .B(N373), .Z(N0) );
  HS65_LH_IVX27 U1152 ( .A(N559), .Z(N1155) );
  HS65_LH_IVX27 U1153 ( .A(N245), .Z(N1152) );
  HS65_LH_AND2X27 U1154 ( .A(N145), .B(N709), .Z(N1147) );
  HS65_LH_IVX49 U1155 ( .A(N2387), .Z(N1141) );
  HS65_LL_AND2X4 U1156 ( .A(N1144), .B(n943), .Z(n509) );
  HS65_LH_OA12X4 U1157 ( .A(n809), .B(n907), .C(n784), .Z(n511) );
  HS65_LL_OR2X9 U1158 ( .A(n1066), .B(n1086), .Z(n522) );
  HS65_LL_MUXI21X2 U1159 ( .D0(n530), .D1(n557), .S0(n556), .Z(n524) );
  HS65_LL_BFX18 U1160 ( .A(N293), .Z(N816) );
  HS65_LH_IVX9 U1161 ( .A(N619), .Z(n874) );
  HS65_LH_MUX21X4 U1162 ( .D0(N341), .D1(N348), .S0(n943), .Z(n948) );
  HS65_LH_IVX9 U1163 ( .A(N523), .Z(n971) );
  HS65_LH_OR2X9 U1164 ( .A(N341), .B(n943), .Z(n528) );
  HS65_LHS_XNOR2X6 U1165 ( .A(n715), .B(n524), .Z(n531) );
  HS65_LH_IVX27 U1166 ( .A(N338), .Z(N1144) );
  HS65_LH_AOI12X6 U1167 ( .A(N348), .B(n943), .C(N523), .Z(n537) );
  HS65_LH_NAND3X2 U1168 ( .A(n952), .B(n637), .C(n753), .Z(n559) );
  HS65_LHS_XNOR2X6 U1169 ( .A(N308), .B(N479), .Z(n573) );
  HS65_LHS_XNOR2X6 U1170 ( .A(N315), .B(N479), .Z(n572) );
  HS65_LH_IVX2 U1171 ( .A(n947), .Z(n575) );
  HS65_LH_NOR2X6 U1172 ( .A(n756), .B(n581), .Z(n673) );
  HS65_LH_IVX9 U1173 ( .A(N625), .Z(n618) );
  HS65_LH_IVX9 U1174 ( .A(N254), .Z(n863) );
  HS65_LH_MUXI21X2 U1175 ( .D0(n863), .D1(n862), .S0(N324), .Z(n601) );
  HS65_LH_MUXI21X2 U1176 ( .D0(N251), .D1(N248), .S0(N324), .Z(n600) );
  HS65_LH_MUXI21X2 U1177 ( .D0(n601), .D1(n600), .S0(N503), .Z(n602) );
  HS65_LH_MUXI21X2 U1178 ( .D0(N251), .D1(N248), .S0(N361), .Z(n977) );
  HS65_LH_IVX9 U1179 ( .A(N248), .Z(n857) );
  HS65_LH_MUXI21X2 U1180 ( .D0(N242), .D1(n857), .S0(N514), .Z(n604) );
  HS65_LH_MUXI21X2 U1181 ( .D0(N254), .D1(N242), .S0(N293), .Z(n999) );
  HS65_LL_MUXI21X2 U1182 ( .D0(N251), .D1(N248), .S0(N302), .Z(n979) );
  HS65_LL_MUXI21X2 U1183 ( .D0(n863), .D1(n862), .S0(N316), .Z(n608) );
  HS65_LL_MUXI21X2 U1184 ( .D0(N251), .D1(N248), .S0(N316), .Z(n607) );
  HS65_LL_MUXI21X2 U1185 ( .D0(n608), .D1(n607), .S0(N490), .Z(n983) );
  HS65_LLS_XOR3X2 U1186 ( .A(n999), .B(n979), .C(n983), .Z(n609) );
  HS65_LH_MUXI21X2 U1187 ( .D0(n863), .D1(n862), .S0(N308), .Z(n613) );
  HS65_LH_MUXI21X2 U1188 ( .D0(N251), .D1(N248), .S0(N308), .Z(n612) );
  HS65_LH_MUXI21X2 U1189 ( .D0(n613), .D1(n612), .S0(N479), .Z(n987) );
  HS65_LHS_XNOR2X6 U1190 ( .A(n614), .B(n987), .Z(n615) );
  HS65_LH_IVX9 U1191 ( .A(N597), .Z(n1007) );
  HS65_LH_IVX9 U1192 ( .A(N598), .Z(n1006) );
  HS65_LH_MUXI41X2 U1193 ( .D0(N596), .D1(n1007), .D2(N595), .D3(n1006), .S0(
        N389), .S1(N257), .Z(n1107) );
  HS65_LH_IVX9 U1194 ( .A(N400), .Z(n801) );
  HS65_LH_OAI21X6 U1195 ( .A(n640), .B(n639), .C(n661), .Z(n754) );
  HS65_LH_MUXI21X2 U1196 ( .D0(N595), .D1(n1006), .S0(N514), .Z(n978) );
  HS65_LH_NOR2X6 U1197 ( .A(N571), .B(n1083), .Z(n645) );
  HS65_LH_NOR2X6 U1198 ( .A(N574), .B(n643), .Z(n1132) );
  HS65_LL_MUXI21X2 U1199 ( .D0(N597), .D1(N598), .S0(N234), .Z(n648) );
  HS65_LH_MUXI31X2 U1200 ( .D0(N596), .D1(N595), .D2(n648), .S0(N234), .S1(
        N435), .Z(n1108) );
  HS65_LH_MUXI21X2 U1201 ( .D0(N257), .D1(N264), .S0(n819), .Z(n653) );
  HS65_LH_MUXI21X2 U1202 ( .D0(N596), .D1(N595), .S0(N324), .Z(n659) );
  HS65_LH_MUXI21X2 U1203 ( .D0(N597), .D1(N598), .S0(N324), .Z(n658) );
  HS65_LL_MX41X14 U1204 ( .D0(n1078), .S0(n1133), .D1(n1079), .S1(n1132), .D2(
        n1131), .S2(N170), .D3(n1130), .S3(N200), .Z(N7600) );
  HS65_LH_NOR2X6 U1205 ( .A(N577), .B(n1083), .Z(n668) );
  HS65_LH_NOR2X6 U1206 ( .A(N580), .B(n666), .Z(n1136) );
  HS65_LH_IVX9 U1207 ( .A(n1117), .Z(n997) );
  HS65_LH_MUX21X9 U1208 ( .D0(N234), .D1(N241), .S0(n819), .Z(n680) );
  HS65_LH_MUXI21X2 U1209 ( .D0(n922), .D1(n921), .S0(N226), .Z(n690) );
  HS65_LH_MUXI21X2 U1210 ( .D0(n690), .D1(n689), .S0(N422), .Z(n1105) );
  HS65_LH_IVX9 U1211 ( .A(N2623), .Z(n1140) );
  HS65_LH_MUXI21X2 U1212 ( .D0(N597), .D1(N598), .S0(N281), .Z(n698) );
  HS65_LH_IVX9 U1213 ( .A(n911), .Z(n699) );
  HS65_LH_NOR2X6 U1214 ( .A(N616), .B(N613), .Z(n1129) );
  HS65_LH_AOI22X4 U1215 ( .A(n762), .B(n995), .C(n1117), .D(n1115), .Z(n721)
         );
  HS65_LL_MUXI21X2 U1216 ( .D0(N596), .D1(N595), .S0(N210), .Z(n726) );
  HS65_LH_IVX9 U1217 ( .A(N457), .Z(n832) );
  HS65_LH_NAND2X7 U1218 ( .A(n730), .B(n832), .Z(n731) );
  HS65_LH_IVX9 U1219 ( .A(n825), .Z(n827) );
  HS65_LH_NAND2X7 U1220 ( .A(n827), .B(n828), .Z(n990) );
  HS65_LH_NAND2X7 U1221 ( .A(n819), .B(n735), .Z(n737) );
  HS65_LH_IVX9 U1222 ( .A(n824), .Z(n839) );
  HS65_LL_OR3ABCX18 U1223 ( .A(n744), .B(n743), .C(n742), .Z(N7740) );
  HS65_LH_NAND4ABX3 U1224 ( .A(n756), .B(n976), .C(n755), .D(n754), .Z(n759)
         );
  HS65_LHS_XNOR2X6 U1225 ( .A(n757), .B(n1116), .Z(n781) );
  HS65_LH_AO12X9 U1226 ( .A(n761), .B(n763), .C(n760), .Z(n998) );
  HS65_LL_AND2X4 U1227 ( .A(n798), .B(n788), .Z(n789) );
  HS65_LHS_XNOR2X6 U1228 ( .A(n796), .B(n815), .Z(n818) );
  HS65_LH_CBI4I1X5 U1229 ( .A(n800), .B(n799), .C(n798), .D(n797), .Z(n814) );
  HS65_LH_MUX21X4 U1230 ( .D0(N273), .D1(N280), .S0(n819), .Z(n935) );
  HS65_LH_MUXI21X2 U1231 ( .D0(n810), .D1(n809), .S0(n905), .Z(n811) );
  HS65_LL_MUXI21X2 U1232 ( .D0(N206), .D1(N209), .S0(n819), .Z(n1017) );
  HS65_LHS_XNOR2X6 U1233 ( .A(n822), .B(n821), .Z(n848) );
  HS65_LH_MUXI21X2 U1234 ( .D0(n1019), .D1(n833), .S0(n839), .Z(n835) );
  HS65_LH_OAI12X3 U1235 ( .A(N619), .B(N118), .C(N625), .Z(n873) );
  HS65_LH_MUXI21X2 U1236 ( .D0(n863), .D1(n862), .S0(N210), .Z(n852) );
  HS65_LH_MUXI21X2 U1237 ( .D0(n852), .D1(n851), .S0(N457), .Z(n854) );
  HS65_LH_MUXI41X2 U1238 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(
        N257), .S1(N389), .Z(n853) );
  HS65_LL_MUXI41X2 U1239 ( .D0(n863), .D1(n862), .D2(N251), .D3(N248), .S0(
        N273), .S1(N411), .Z(n859) );
  HS65_LH_MUXI21X2 U1240 ( .D0(N596), .D1(N595), .S0(N218), .Z(n883) );
  HS65_LH_MUXI21X2 U1241 ( .D0(N597), .D1(N598), .S0(N218), .Z(n881) );
  HS65_LH_OAI21X3 U1242 ( .A(N468), .B(n883), .C(n882), .Z(n1104) );
  HS65_LH_IVX9 U1243 ( .A(n885), .Z(n889) );
  HS65_LH_NAND2X7 U1244 ( .A(n1128), .B(n1075), .Z(n896) );
  HS65_LH_NOR4ABX2 U1245 ( .A(n926), .B(n911), .C(n1009), .D(n910), .Z(n912)
         );
  HS65_LL_AND3ABCX18 U1246 ( .A(n920), .B(n919), .C(n1003), .Z(N7503) );
  HS65_LH_MUXI21X2 U1247 ( .D0(n922), .D1(n921), .S0(N273), .Z(n924) );
  HS65_LH_MUXI21X2 U1248 ( .D0(N597), .D1(N598), .S0(N273), .Z(n923) );
  HS65_LH_MUXI21X2 U1249 ( .D0(n924), .D1(n923), .S0(N411), .Z(n1110) );
  HS65_LHS_XOR3X2 U1250 ( .A(n931), .B(n930), .C(n929), .Z(n942) );
  HS65_LH_MUXI21X2 U1251 ( .D0(n961), .D1(n938), .S0(n937), .Z(n939) );
  HS65_LL_XNOR2X18 U1252 ( .A(n942), .B(n941), .Z(N7476) );
  HS65_LH_BFX49 U1253 ( .A(N299), .Z(N2527) );
  HS65_LH_MUXI21X2 U1254 ( .D0(n945), .D1(n944), .S0(n943), .Z(n946) );
  HS65_LHS_XOR3X2 U1255 ( .A(n948), .B(n947), .C(n946), .Z(n955) );
  HS65_LH_MUXI21X2 U1256 ( .D0(n950), .D1(N331), .S0(n949), .Z(n951) );
  HS65_LHS_XOR3X2 U1257 ( .A(n953), .B(n952), .C(n951), .Z(n954) );
  HS65_LHS_XNOR3X2 U1258 ( .A(n962), .B(n961), .C(n960), .Z(n963) );
  HS65_LHS_XOR3X2 U1259 ( .A(N324), .B(N316), .C(n965), .Z(n968) );
  HS65_LHS_XOR3X2 U1260 ( .A(N369), .B(N361), .C(N816), .Z(n966) );
  HS65_LHS_XOR3X2 U1261 ( .A(N302), .B(N308), .C(n966), .Z(n967) );
  HS65_LL_NAND4ABX3 U1262 ( .A(N6877), .B(n1094), .C(N1140), .D(n969), .Z(n970) );
  HS65_LL_AND3ABCX18 U1263 ( .A(N7474), .B(n970), .C(N7476), .Z(N7703) );
  HS65_LH_MUXI21X2 U1264 ( .D0(n1007), .D1(n1006), .S0(N341), .Z(n973) );
  HS65_LH_MUXI21X2 U1265 ( .D0(N596), .D1(N595), .S0(N341), .Z(n972) );
  HS65_LH_MUXI21X2 U1266 ( .D0(n973), .D1(n972), .S0(n971), .Z(n982) );
  HS65_LH_NOR4ABX2 U1267 ( .A(n999), .B(n980), .C(n979), .D(n978), .Z(n981) );
  HS65_LL_AND2ABX27 U1268 ( .A(n993), .B(n1022), .Z(N6648) );
  HS65_LL_AO112X27 U1269 ( .A(n997), .B(n996), .C(n995), .D(n994), .Z(N6927)
         );
  HS65_LL_MX41X14 U1270 ( .D0(n1122), .S0(n1129), .D1(n1121), .S1(n1128), .D2(
        n711), .S2(N106), .D3(n1127), .S3(N109), .Z(N7735) );
  HS65_LL_MX41X14 U1271 ( .D0(n1114), .S0(n1129), .D1(n1060), .S1(n1128), .D2(
        n711), .S2(N40), .D3(n1127), .S3(N91), .Z(N7742) );
  HS65_LL_MX41X14 U1272 ( .D0(n1030), .S0(n1129), .D1(n1064), .S1(n1128), .D2(
        n711), .S2(N20), .D3(n1127), .S3(N76), .Z(N7520) );
  HS65_LL_MX41X14 U1273 ( .D0(n1079), .S0(n1129), .D1(n1078), .S1(n1128), .D2(
        n711), .S2(N37), .D3(n1127), .S3(N43), .Z(N7519) );
  HS65_LL_AND2ABX18 U1274 ( .A(n1016), .B(n519), .Z(N7472) );
  HS65_LH_NOR2X6 U1275 ( .A(N607), .B(N610), .Z(n1126) );
  HS65_LH_NOR2X6 U1276 ( .A(N607), .B(n1028), .Z(n1125) );
  HS65_LH_IVX71 U1277 ( .A(N545), .Z(N1137) );
  HS65_LL_NAND2X14 U1278 ( .A(n1047), .B(n1046), .Z(N8124) );
  HS65_LH_MUXI21X2 U1279 ( .D0(N176), .D1(N179), .S0(N577), .Z(n1067) );
  HS65_LH_MUXI21X2 U1280 ( .D0(N176), .D1(N179), .S0(N571), .Z(n1084) );
  HS65_LH_MUXI21X2 U1281 ( .D0(n1098), .D1(N123), .S0(N599), .Z(n1099) );
  HS65_LH_OR4X4 U1282 ( .A(n1110), .B(n1109), .C(n1108), .D(n1107), .Z(n1111)
         );
  HS65_LL_MX41X14 U1283 ( .D0(n508), .S0(n1129), .D1(n1123), .S1(n1128), .D2(
        n711), .S2(N70), .D3(n1127), .S3(N67), .Z(N7522) );
  HS65_LL_MX41X14 U1284 ( .D0(n700), .S0(n1133), .D1(n507), .S1(n1132), .D2(
        n1131), .S2(N185), .D3(n1130), .S3(N182), .Z(N7506) );
  HS65_LL_MX41X14 U1285 ( .D0(n700), .S0(n1138), .D1(n507), .S1(n1136), .D2(
        n1135), .S2(N185), .D3(n1134), .S3(N182), .Z(N7511) );
  HS65_LL_MX41X14 U1286 ( .D0(n507), .S0(n1126), .D1(n700), .S1(n1125), .D2(
        n1029), .S2(N61), .D3(n1124), .S3(N11), .Z(N7449) );
  HS65_LL_MX41X14 U1287 ( .D0(n507), .S0(n1129), .D1(n700), .S1(n1128), .D2(
        n711), .S2(N61), .D3(n1127), .S3(N11), .Z(N7469) );
  HS65_LL_MX41X14 U1288 ( .D0(n1123), .S0(n1133), .D1(n508), .S1(n1132), .D2(
        n1131), .S2(N158), .D3(n1130), .S3(N188), .Z(N7601) );
  HS65_LL_MX41X14 U1289 ( .D0(n1123), .S0(n1138), .D1(n508), .S1(n1136), .D2(
        n1135), .S2(N158), .D3(n1134), .S3(N188), .Z(N7605) );
  HS65_LL_MX41X14 U1290 ( .D0(n1137), .S0(n1126), .D1(n1139), .S1(n1125), .D2(
        n1029), .S2(N17), .D3(n1124), .S3(N73), .Z(N7517) );
  HS65_LL_MX41X14 U1291 ( .D0(n1137), .S0(n1129), .D1(n1139), .S1(n1128), .D2(
        n711), .S2(N17), .D3(n1127), .S3(N73), .Z(N7521) );
  HS65_LL_MX41X14 U1292 ( .D0(n1139), .S0(n1133), .D1(n1137), .S1(n1132), .D2(
        n1131), .S2(N152), .D3(n1130), .S3(N155), .Z(N7602) );
  HS65_LL_MX41X14 U1293 ( .D0(n1139), .S0(n1138), .D1(n1137), .S1(n1136), .D2(
        n1135), .S2(N152), .D3(n1134), .S3(N155), .Z(N7606) );
endmodule

