
module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   N0, N23, N34, N35, N36, N37, N38, N39, N40, N41, N50, N51, N52, N53,
         N54, N55, N56, N57, N66, N67, N68, N69, N70, N71, N72, N73, N82, N83,
         N84, N85, N86, N87, N88, N89, N98, N99, N100, N101, N102, N103, N104,
         N105, N114, N115, N116, N117, N118, N119, N120, N121, N130, N131,
         N132, N133, N134, N135, N136, N137, N146, N147, N148, N149, N150,
         N151, N152, N153, N162, N163, N164, N165, N166, N167, N168, N169,
         N178, N179, N180, N181, N182, N183, N184, N185, N194, N195, N196,
         N197, N198, N199, N200, N201, N210, N211, N212, N213, N214, N215,
         N216, N217, N226, N227, N228, N229, N230, N231, N232, N233, N242,
         N243, N244, N245, N246, N247, N248, N249, N258, N259, N260, N261,
         N262, N263, N264, N265, N274, N275, N276, N277, N278, N279, N280,
         N281, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, \u0/N271 , \u0/N270 ,
         \u0/N269 , \u0/N268 , \u0/N267 , \u0/N266 , \u0/N265 , \u0/N264 ,
         \u0/N263 , \u0/N262 , \u0/N261 , \u0/N260 , \u0/N259 , \u0/N258 ,
         \u0/N257 , \u0/N256 , \u0/N255 , \u0/N254 , \u0/N253 , \u0/N252 ,
         \u0/N251 , \u0/N250 , \u0/N249 , \u0/N248 , \u0/N247 , \u0/N246 ,
         \u0/N245 , \u0/N244 , \u0/N243 , \u0/N242 , \u0/N241 , \u0/N240 ,
         \u0/N205 , \u0/N204 , \u0/N203 , \u0/N202 , \u0/N201 , \u0/N200 ,
         \u0/N199 , \u0/N198 , \u0/N197 , \u0/N196 , \u0/N195 , \u0/N194 ,
         \u0/N193 , \u0/N192 , \u0/N191 , \u0/N190 , \u0/N189 , \u0/N188 ,
         \u0/N187 , \u0/N186 , \u0/N185 , \u0/N184 , \u0/N183 , \u0/N182 ,
         \u0/N181 , \u0/N180 , \u0/N179 , \u0/N178 , \u0/N177 , \u0/N176 ,
         \u0/N175 , \u0/N174 , \u0/N139 , \u0/N138 , \u0/N137 , \u0/N136 ,
         \u0/N135 , \u0/N134 , \u0/N133 , \u0/N132 , \u0/N131 , \u0/N130 ,
         \u0/N129 , \u0/N128 , \u0/N127 , \u0/N126 , \u0/N125 , \u0/N124 ,
         \u0/N123 , \u0/N122 , \u0/N121 , \u0/N120 , \u0/N119 , \u0/N118 ,
         \u0/N117 , \u0/N116 , \u0/N115 , \u0/N114 , \u0/N113 , \u0/N112 ,
         \u0/N111 , \u0/N110 , \u0/N109 , \u0/N108 , \u0/N73 , \u0/N72 ,
         \u0/N71 , \u0/N70 , \u0/N69 , \u0/N68 , \u0/N67 , \u0/N66 , \u0/N65 ,
         \u0/N64 , \u0/N63 , \u0/N62 , \u0/N61 , \u0/N60 , \u0/N59 , \u0/N58 ,
         \u0/N57 , \u0/N56 , \u0/N55 , \u0/N54 , \u0/N53 , \u0/N52 , \u0/N51 ,
         \u0/N50 , \u0/N49 , \u0/N48 , \u0/N47 , \u0/N46 , \u0/N45 , \u0/N44 ,
         \u0/N43 , \u0/N42 , \u0/r0/N81 , \u0/r0/N80 , \u0/r0/N79 ,
         \u0/r0/N78 , \u0/r0/N77 , \u0/r0/N76 , \u0/r0/N75 , \u0/r0/N74 ,
         \u0/r0/N73 , \u0/r0/N72 , \u0/r0/N71 , \u0/r0/N70 , n1, n2, n3, n4,
         n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n928, n930, n931, n933, n934, n938,
         n939, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa23;
  wire   [7:0] sa13;
  wire   [7:0] sa03;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa22;
  wire   [7:0] sa12;
  wire   [7:0] sa02;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa21;
  wire   [7:0] sa11;
  wire   [7:0] sa01;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa20;
  wire   [7:0] sa10;
  wire   [7:0] sa00;
  wire   [31:0] \u0/rcon ;
  wire   [3:0] \u0/r0/rcnt ;

  HS65_LL_DFPQX4 \dcnt_reg[0]  ( .D(n9114), .CP(clk), .Q(dcnt[0]) );
  HS65_LL_DFPQX4 \dcnt_reg[1]  ( .D(n9112), .CP(clk), .Q(dcnt[1]) );
  HS65_LL_DFPQX4 \dcnt_reg[2]  ( .D(n9111), .CP(clk), .Q(dcnt[2]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[0]  ( .D(\u0/r0/N78 ), .CP(clk), .Q(
        \u0/r0/rcnt [0]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[1]  ( .D(\u0/r0/N79 ), .CP(clk), .Q(
        \u0/r0/rcnt [1]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[2]  ( .D(\u0/r0/N80 ), .CP(clk), .Q(
        \u0/r0/rcnt [2]) );
  HS65_LL_DFPQX4 \u0/r0/rcnt_reg[3]  ( .D(\u0/r0/N81 ), .CP(clk), .Q(
        \u0/r0/rcnt [3]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[24]  ( .D(\u0/r0/N70 ), .CP(clk), .Q(
        \u0/rcon [24]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[25]  ( .D(\u0/r0/N71 ), .CP(clk), .Q(
        \u0/rcon [25]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[26]  ( .D(\u0/r0/N72 ), .CP(clk), .Q(
        \u0/rcon [26]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[27]  ( .D(\u0/r0/N73 ), .CP(clk), .Q(
        \u0/rcon [27]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[28]  ( .D(\u0/r0/N74 ), .CP(clk), .Q(
        \u0/rcon [28]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[29]  ( .D(\u0/r0/N75 ), .CP(clk), .Q(
        \u0/rcon [29]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[30]  ( .D(\u0/r0/N76 ), .CP(clk), .Q(
        \u0/rcon [30]) );
  HS65_LL_DFPQX4 \u0/r0/out_reg[31]  ( .D(\u0/r0/N77 ), .CP(clk), .Q(
        \u0/rcon [31]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][31]  ( .D(\u0/N73 ), .CP(clk), .Q(w0[31]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][31]  ( .D(\u0/N271 ), .CP(clk), .Q(w3[31]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][0]  ( .D(\u0/N42 ), .CP(clk), .Q(w0[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][0]  ( .D(\u0/N240 ), .CP(clk), .Q(w3[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][8]  ( .D(\u0/N50 ), .CP(clk), .Q(w0[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][8]  ( .D(\u0/N248 ), .CP(clk), .Q(w3[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][16]  ( .D(\u0/N58 ), .CP(clk), .Q(w0[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][16]  ( .D(\u0/N256 ), .CP(clk), .Q(w3[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][24]  ( .D(\u0/N66 ), .CP(clk), .Q(w0[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][24]  ( .D(\u0/N264 ), .CP(clk), .Q(w3[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][3]  ( .D(\u0/N45 ), .CP(clk), .Q(w0[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][3]  ( .D(\u0/N243 ), .CP(clk), .Q(w3[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][10]  ( .D(\u0/N52 ), .CP(clk), .Q(w0[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][10]  ( .D(\u0/N250 ), .CP(clk), .Q(w3[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][23]  ( .D(\u0/N65 ), .CP(clk), .Q(w0[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][23]  ( .D(\u0/N263 ), .CP(clk), .Q(w3[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][25]  ( .D(\u0/N67 ), .CP(clk), .Q(w0[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][25]  ( .D(\u0/N265 ), .CP(clk), .Q(w3[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][7]  ( .D(\u0/N49 ), .CP(clk), .Q(w0[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][7]  ( .D(\u0/N247 ), .CP(clk), .Q(w3[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][9]  ( .D(\u0/N51 ), .CP(clk), .Q(w0[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][9]  ( .D(\u0/N249 ), .CP(clk), .Q(w3[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][18]  ( .D(\u0/N60 ), .CP(clk), .Q(w0[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][18]  ( .D(\u0/N258 ), .CP(clk), .Q(w3[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][27]  ( .D(\u0/N69 ), .CP(clk), .Q(w0[27]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][27]  ( .D(\u0/N267 ), .CP(clk), .Q(w3[27]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][2]  ( .D(\u0/N44 ), .CP(clk), .Q(w0[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][2]  ( .D(\u0/N242 ), .CP(clk), .Q(w3[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][15]  ( .D(\u0/N57 ), .CP(clk), .Q(w0[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][15]  ( .D(\u0/N255 ), .CP(clk), .Q(w3[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][17]  ( .D(\u0/N59 ), .CP(clk), .Q(w0[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][17]  ( .D(\u0/N257 ), .CP(clk), .Q(w3[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][26]  ( .D(\u0/N68 ), .CP(clk), .Q(w0[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][26]  ( .D(\u0/N266 ), .CP(clk), .Q(w3[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][6]  ( .D(\u0/N48 ), .CP(clk), .Q(w0[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][6]  ( .D(\u0/N246 ), .CP(clk), .Q(w3[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][11]  ( .D(\u0/N53 ), .CP(clk), .Q(w0[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][11]  ( .D(\u0/N251 ), .CP(clk), .Q(w3[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][19]  ( .D(\u0/N61 ), .CP(clk), .Q(w0[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][19]  ( .D(\u0/N259 ), .CP(clk), .Q(w3[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][30]  ( .D(\u0/N72 ), .CP(clk), .Q(w0[30]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][30]  ( .D(\u0/N270 ), .CP(clk), .Q(w3[30]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][4]  ( .D(\u0/N46 ), .CP(clk), .Q(w0[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][4]  ( .D(\u0/N244 ), .CP(clk), .Q(w3[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][13]  ( .D(\u0/N55 ), .CP(clk), .Q(w0[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][13]  ( .D(\u0/N253 ), .CP(clk), .Q(w3[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][21]  ( .D(\u0/N63 ), .CP(clk), .Q(w0[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][21]  ( .D(\u0/N261 ), .CP(clk), .Q(w3[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][29]  ( .D(\u0/N71 ), .CP(clk), .Q(w0[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][29]  ( .D(\u0/N269 ), .CP(clk), .Q(w3[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][5]  ( .D(\u0/N47 ), .CP(clk), .Q(w0[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][5]  ( .D(\u0/N245 ), .CP(clk), .Q(w3[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][12]  ( .D(\u0/N54 ), .CP(clk), .Q(w0[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][12]  ( .D(\u0/N252 ), .CP(clk), .Q(w3[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][22]  ( .D(\u0/N64 ), .CP(clk), .Q(w0[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][22]  ( .D(\u0/N262 ), .CP(clk), .Q(w3[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][28]  ( .D(\u0/N70 ), .CP(clk), .Q(w0[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][28]  ( .D(\u0/N268 ), .CP(clk), .Q(w3[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][1]  ( .D(\u0/N43 ), .CP(clk), .Q(w0[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][1]  ( .D(\u0/N241 ), .CP(clk), .Q(w3[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][14]  ( .D(\u0/N56 ), .CP(clk), .Q(w0[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][14]  ( .D(\u0/N254 ), .CP(clk), .Q(w3[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[0][20]  ( .D(\u0/N62 ), .CP(clk), .Q(w0[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[3][20]  ( .D(\u0/N260 ), .CP(clk), .Q(w3[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][20]  ( .D(\u0/N194 ), .CP(clk), .Q(w2[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][20]  ( .D(\u0/N128 ), .CP(clk), .Q(w1[20]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][14]  ( .D(\u0/N188 ), .CP(clk), .Q(w2[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][14]  ( .D(\u0/N122 ), .CP(clk), .Q(w1[14]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][1]  ( .D(\u0/N175 ), .CP(clk), .Q(w2[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][1]  ( .D(\u0/N109 ), .CP(clk), .Q(w1[1]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][28]  ( .D(\u0/N202 ), .CP(clk), .Q(w2[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][28]  ( .D(\u0/N136 ), .CP(clk), .Q(w1[28]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][22]  ( .D(\u0/N196 ), .CP(clk), .Q(w2[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][22]  ( .D(\u0/N130 ), .CP(clk), .Q(w1[22]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][12]  ( .D(\u0/N186 ), .CP(clk), .Q(w2[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][12]  ( .D(\u0/N120 ), .CP(clk), .Q(w1[12]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][5]  ( .D(\u0/N179 ), .CP(clk), .Q(w2[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][5]  ( .D(\u0/N113 ), .CP(clk), .Q(w1[5]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][29]  ( .D(\u0/N203 ), .CP(clk), .Q(w2[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][29]  ( .D(\u0/N137 ), .CP(clk), .Q(w1[29]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][21]  ( .D(\u0/N195 ), .CP(clk), .Q(w2[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][21]  ( .D(\u0/N129 ), .CP(clk), .Q(w1[21]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][13]  ( .D(\u0/N187 ), .CP(clk), .Q(w2[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][13]  ( .D(\u0/N121 ), .CP(clk), .Q(w1[13]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][4]  ( .D(\u0/N178 ), .CP(clk), .Q(w2[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][4]  ( .D(\u0/N112 ), .CP(clk), .Q(w1[4]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][30]  ( .D(\u0/N204 ), .CP(clk), .Q(w2[30]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][30]  ( .D(\u0/N138 ), .CP(clk), .Q(w1[30]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][19]  ( .D(\u0/N193 ), .CP(clk), .Q(w2[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][19]  ( .D(\u0/N127 ), .CP(clk), .Q(w1[19]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][11]  ( .D(\u0/N185 ), .CP(clk), .Q(w2[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][11]  ( .D(\u0/N119 ), .CP(clk), .Q(w1[11]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][6]  ( .D(\u0/N180 ), .CP(clk), .Q(w2[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][6]  ( .D(\u0/N114 ), .CP(clk), .Q(w1[6]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][26]  ( .D(\u0/N200 ), .CP(clk), .Q(w2[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][26]  ( .D(\u0/N134 ), .CP(clk), .Q(w1[26]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][17]  ( .D(\u0/N191 ), .CP(clk), .Q(w2[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][17]  ( .D(\u0/N125 ), .CP(clk), .Q(w1[17]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][15]  ( .D(\u0/N189 ), .CP(clk), .Q(w2[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][15]  ( .D(\u0/N123 ), .CP(clk), .Q(w1[15]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][2]  ( .D(\u0/N176 ), .CP(clk), .Q(w2[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][2]  ( .D(\u0/N110 ), .CP(clk), .Q(w1[2]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][27]  ( .D(\u0/N201 ), .CP(clk), .Q(w2[27]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][27]  ( .D(\u0/N135 ), .CP(clk), .Q(w1[27]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][18]  ( .D(\u0/N192 ), .CP(clk), .Q(w2[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][18]  ( .D(\u0/N126 ), .CP(clk), .Q(w1[18]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][9]  ( .D(\u0/N183 ), .CP(clk), .Q(w2[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][9]  ( .D(\u0/N117 ), .CP(clk), .Q(w1[9]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][7]  ( .D(\u0/N181 ), .CP(clk), .Q(w2[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][7]  ( .D(\u0/N115 ), .CP(clk), .Q(w1[7]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][25]  ( .D(\u0/N199 ), .CP(clk), .Q(w2[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][25]  ( .D(\u0/N133 ), .CP(clk), .Q(w1[25]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][23]  ( .D(\u0/N197 ), .CP(clk), .Q(w2[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][23]  ( .D(\u0/N131 ), .CP(clk), .Q(w1[23]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][10]  ( .D(\u0/N184 ), .CP(clk), .Q(w2[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][10]  ( .D(\u0/N118 ), .CP(clk), .Q(w1[10]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][3]  ( .D(\u0/N177 ), .CP(clk), .Q(w2[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][3]  ( .D(\u0/N111 ), .CP(clk), .Q(w1[3]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][24]  ( .D(\u0/N198 ), .CP(clk), .Q(w2[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][24]  ( .D(\u0/N132 ), .CP(clk), .Q(w1[24]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][16]  ( .D(\u0/N190 ), .CP(clk), .Q(w2[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][16]  ( .D(\u0/N124 ), .CP(clk), .Q(w1[16]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][8]  ( .D(\u0/N182 ), .CP(clk), .Q(w2[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][8]  ( .D(\u0/N116 ), .CP(clk), .Q(w1[8]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][0]  ( .D(\u0/N174 ), .CP(clk), .Q(w2[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][0]  ( .D(\u0/N108 ), .CP(clk), .Q(w1[0]) );
  HS65_LL_DFPQX4 \u0/w_reg[2][31]  ( .D(\u0/N205 ), .CP(clk), .Q(w2[31]) );
  HS65_LL_DFPQX4 \u0/w_reg[1][31]  ( .D(\u0/N139 ), .CP(clk), .Q(w1[31]) );
  HS65_LL_DFPQX4 \sa01_reg[7]  ( .D(N217), .CP(clk), .Q(sa01[7]) );
  HS65_LL_DFPQX4 \sa31_reg[0]  ( .D(N162), .CP(clk), .Q(sa31[0]) );
  HS65_LL_DFPQX4 \sa32_reg[2]  ( .D(N100), .CP(clk), .Q(sa32[2]) );
  HS65_LL_DFPQX4 \sa33_reg[0]  ( .D(N34), .CP(clk), .Q(sa33[0]) );
  HS65_LL_DFPQX4 \sa30_reg[0]  ( .D(N226), .CP(clk), .Q(sa30[0]) );
  HS65_LL_DFPQX4 \sa21_reg[3]  ( .D(N181), .CP(clk), .Q(sa21[3]) );
  HS65_LL_DFPQX4 \sa13_reg[1]  ( .D(N67), .CP(clk), .Q(sa13[1]) );
  HS65_LL_DFPQX4 \sa12_reg[3]  ( .D(N133), .CP(clk), .Q(sa12[3]) );
  HS65_LL_DFPQX4 \sa11_reg[1]  ( .D(N195), .CP(clk), .Q(sa11[1]) );
  HS65_LL_DFPQX4 \sa10_reg[1]  ( .D(N259), .CP(clk), .Q(sa10[1]) );
  HS65_LL_DFPQX4 \sa23_reg[0]  ( .D(N50), .CP(clk), .Q(sa23[0]) );
  HS65_LL_DFPQX4 \sa21_reg[1]  ( .D(N179), .CP(clk), .Q(sa21[1]) );
  HS65_LL_DFPQX4 \sa23_reg[1]  ( .D(N51), .CP(clk), .Q(sa23[1]) );
  HS65_LL_DFPQX4 \sa31_reg[2]  ( .D(N164), .CP(clk), .Q(sa31[2]) );
  HS65_LL_DFPQX4 \sa32_reg[3]  ( .D(N101), .CP(clk), .Q(sa32[3]) );
  HS65_LL_DFPQX4 \sa33_reg[3]  ( .D(N37), .CP(clk), .Q(sa33[3]) );
  HS65_LL_DFPQX4 \sa30_reg[4]  ( .D(N230), .CP(clk), .Q(sa30[4]) );
  HS65_LL_DFPQX4 \sa31_reg[3]  ( .D(N165), .CP(clk), .Q(sa31[3]) );
  HS65_LL_DFPQX4 \sa12_reg[2]  ( .D(N132), .CP(clk), .Q(sa12[2]) );
  HS65_LL_DFPQX4 \sa11_reg[0]  ( .D(N194), .CP(clk), .Q(sa11[0]) );
  HS65_LL_DFPQX4 \sa30_reg[3]  ( .D(N229), .CP(clk), .Q(sa30[3]) );
  HS65_LL_DFPQX4 \sa31_reg[4]  ( .D(N166), .CP(clk), .Q(sa31[4]) );
  HS65_LL_DFPQX4 \sa22_reg[0]  ( .D(N114), .CP(clk), .Q(sa22[0]) );
  HS65_LL_DFPQX4 \sa20_reg[1]  ( .D(N243), .CP(clk), .Q(sa20[1]) );
  HS65_LL_DFPQX4 \sa22_reg[3]  ( .D(N117), .CP(clk), .Q(sa22[3]) );
  HS65_LL_DFPQX4 \sa30_reg[1]  ( .D(N227), .CP(clk), .Q(sa30[1]) );
  HS65_LL_DFPQX4 \sa01_reg[0]  ( .D(N210), .CP(clk), .Q(sa01[0]) );
  HS65_LL_DFPQX4 \sa21_reg[0]  ( .D(N178), .CP(clk), .Q(sa21[0]) );
  HS65_LL_DFPQX4 \sa31_reg[1]  ( .D(N163), .CP(clk), .Q(sa31[1]) );
  HS65_LL_DFPQX4 \sa22_reg[4]  ( .D(N118), .CP(clk), .Q(sa22[4]) );
  HS65_LL_DFPQX4 \sa30_reg[7]  ( .D(N233), .CP(clk), .Q(sa30[7]) );
  HS65_LL_DFPQX4 \sa31_reg[5]  ( .D(N167), .CP(clk), .Q(sa31[5]) );
  HS65_LL_DFPQX4 \sa32_reg[7]  ( .D(N105), .CP(clk), .Q(sa32[7]) );
  HS65_LL_DFPQX4 \sa03_reg[4]  ( .D(N86), .CP(clk), .Q(sa03[4]) );
  HS65_LL_DFPQX4 \sa33_reg[7]  ( .D(N41), .CP(clk), .Q(sa33[7]) );
  HS65_LL_DFPQX4 \sa30_reg[5]  ( .D(N231), .CP(clk), .Q(sa30[5]) );
  HS65_LL_DFPQX4 \sa31_reg[7]  ( .D(N169), .CP(clk), .Q(sa31[7]) );
  HS65_LL_DFPQX4 \sa32_reg[5]  ( .D(N103), .CP(clk), .Q(sa32[5]) );
  HS65_LL_DFPQX4 \sa33_reg[4]  ( .D(N38), .CP(clk), .Q(sa33[4]) );
  HS65_LL_DFPQX4 \sa20_reg[2]  ( .D(N244), .CP(clk), .Q(sa20[2]) );
  HS65_LL_DFPQX4 \sa22_reg[2]  ( .D(N116), .CP(clk), .Q(sa22[2]) );
  HS65_LL_DFPQX4 \sa12_reg[1]  ( .D(N131), .CP(clk), .Q(sa12[1]) );
  HS65_LL_DFPQX4 \sa11_reg[2]  ( .D(N196), .CP(clk), .Q(sa11[2]) );
  HS65_LL_DFPQX4 \sa30_reg[2]  ( .D(N228), .CP(clk), .Q(sa30[2]) );
  HS65_LL_DFPQX4 \sa31_reg[6]  ( .D(N168), .CP(clk), .Q(sa31[6]) );
  HS65_LL_DFPQX4 \sa22_reg[6]  ( .D(N120), .CP(clk), .Q(sa22[6]) );
  HS65_LL_DFPQX4 \sa10_reg[2]  ( .D(N260), .CP(clk), .Q(sa10[2]) );
  HS65_LL_DFPQX4 \sa20_reg[3]  ( .D(N245), .CP(clk), .Q(sa20[3]) );
  HS65_LL_DFPQX4 \sa22_reg[1]  ( .D(N115), .CP(clk), .Q(sa22[1]) );
  HS65_LL_DFPQX4 \sa10_reg[5]  ( .D(N263), .CP(clk), .Q(sa10[5]) );
  HS65_LL_DFPQX4 \sa03_reg[2]  ( .D(N84), .CP(clk), .Q(sa03[2]) );
  HS65_LL_DFPQX4 \sa33_reg[1]  ( .D(N35), .CP(clk), .Q(sa33[1]) );
  HS65_LL_DFPQX4 \sa20_reg[0]  ( .D(N242), .CP(clk), .Q(sa20[0]) );
  HS65_LL_DFPQX4 \sa12_reg[0]  ( .D(N130), .CP(clk), .Q(sa12[0]) );
  HS65_LL_DFPQX4 \sa11_reg[4]  ( .D(N198), .CP(clk), .Q(sa11[4]) );
  HS65_LL_DFPQX4 \sa10_reg[6]  ( .D(N264), .CP(clk), .Q(sa10[6]) );
  HS65_LL_DFPQX4 \sa23_reg[2]  ( .D(N52), .CP(clk), .Q(sa23[2]) );
  HS65_LL_DFPQX4 \sa21_reg[2]  ( .D(N180), .CP(clk), .Q(sa21[2]) );
  HS65_LL_DFPQX4 \sa13_reg[4]  ( .D(N70), .CP(clk), .Q(sa13[4]) );
  HS65_LL_DFPQX4 \sa02_reg[1]  ( .D(N147), .CP(clk), .Q(sa02[1]) );
  HS65_LL_DFPQX4 \sa32_reg[1]  ( .D(N99), .CP(clk), .Q(sa32[1]) );
  HS65_LL_DFPQX4 \sa02_reg[2]  ( .D(N148), .CP(clk), .Q(sa02[2]) );
  HS65_LL_DFPQX4 \sa02_reg[3]  ( .D(N149), .CP(clk), .Q(sa02[3]) );
  HS65_LL_DFPQX4 \sa32_reg[6]  ( .D(N104), .CP(clk), .Q(sa32[6]) );
  HS65_LL_DFPQX4 \sa23_reg[7]  ( .D(N57), .CP(clk), .Q(sa23[7]) );
  HS65_LL_DFPQX4 \sa11_reg[5]  ( .D(N199), .CP(clk), .Q(sa11[5]) );
  HS65_LL_DFPQX4 \sa10_reg[4]  ( .D(N262), .CP(clk), .Q(sa10[4]) );
  HS65_LL_DFPQX4 \sa10_reg[0]  ( .D(N258), .CP(clk), .Q(sa10[0]) );
  HS65_LL_DFPQX4 \sa13_reg[0]  ( .D(N66), .CP(clk), .Q(sa13[0]) );
  HS65_LL_DFPQX4 \sa02_reg[0]  ( .D(N146), .CP(clk), .Q(sa02[0]) );
  HS65_LL_DFPQX4 \sa32_reg[0]  ( .D(N98), .CP(clk), .Q(sa32[0]) );
  HS65_LL_DFPQX4 \sa03_reg[0]  ( .D(N82), .CP(clk), .Q(sa03[0]) );
  HS65_LL_DFPQX4 \sa03_reg[3]  ( .D(N85), .CP(clk), .Q(sa03[3]) );
  HS65_LL_DFPQX4 \sa33_reg[2]  ( .D(N36), .CP(clk), .Q(sa33[2]) );
  HS65_LL_DFPQX4 \sa20_reg[5]  ( .D(N247), .CP(clk), .Q(sa20[5]) );
  HS65_LL_DFPQX4 \sa12_reg[6]  ( .D(N136), .CP(clk), .Q(sa12[6]) );
  HS65_LL_DFPQX4 \sa21_reg[5]  ( .D(N183), .CP(clk), .Q(sa21[5]) );
  HS65_LL_DFPQX4 \sa11_reg[6]  ( .D(N200), .CP(clk), .Q(sa11[6]) );
  HS65_LL_DFPQX4 \sa20_reg[4]  ( .D(N246), .CP(clk), .Q(sa20[4]) );
  HS65_LL_DFPQX4 \sa12_reg[5]  ( .D(N135), .CP(clk), .Q(sa12[5]) );
  HS65_LL_DFPQX4 \sa32_reg[4]  ( .D(N102), .CP(clk), .Q(sa32[4]) );
  HS65_LL_DFPQX4 \sa03_reg[1]  ( .D(N83), .CP(clk), .Q(sa03[1]) );
  HS65_LL_DFPQX4 \sa33_reg[5]  ( .D(N39), .CP(clk), .Q(sa33[5]) );
  HS65_LL_DFPQX4 \sa20_reg[6]  ( .D(N248), .CP(clk), .Q(sa20[6]) );
  HS65_LL_DFPQX4 \sa12_reg[4]  ( .D(N134), .CP(clk), .Q(sa12[4]) );
  HS65_LL_DFPQX4 \sa21_reg[4]  ( .D(N182), .CP(clk), .Q(sa21[4]) );
  HS65_LL_DFPQX4 \sa13_reg[2]  ( .D(N68), .CP(clk), .Q(sa13[2]) );
  HS65_LL_DFPQX4 \sa02_reg[4]  ( .D(N150), .CP(clk), .Q(sa02[4]) );
  HS65_LL_DFPQX4 \sa22_reg[7]  ( .D(N121), .CP(clk), .Q(sa22[7]) );
  HS65_LL_DFPQX4 \sa10_reg[3]  ( .D(N261), .CP(clk), .Q(sa10[3]) );
  HS65_LL_DFPQX4 \sa23_reg[4]  ( .D(N54), .CP(clk), .Q(sa23[4]) );
  HS65_LL_DFPQX4 \sa13_reg[5]  ( .D(N71), .CP(clk), .Q(sa13[5]) );
  HS65_LL_DFPQX4 \sa12_reg[7]  ( .D(N137), .CP(clk), .Q(sa12[7]) );
  HS65_LL_DFPQX4 \sa11_reg[7]  ( .D(N201), .CP(clk), .Q(sa11[7]) );
  HS65_LL_DFPQX4 \sa00_reg[2]  ( .D(N276), .CP(clk), .Q(sa00[2]) );
  HS65_LL_DFPQX4 \sa10_reg[7]  ( .D(N265), .CP(clk), .Q(sa10[7]) );
  HS65_LL_DFPQX4 \sa23_reg[5]  ( .D(N55), .CP(clk), .Q(sa23[5]) );
  HS65_LL_DFPQX4 \sa21_reg[7]  ( .D(N185), .CP(clk), .Q(sa21[7]) );
  HS65_LL_DFPQX4 \sa23_reg[3]  ( .D(N53), .CP(clk), .Q(sa23[3]) );
  HS65_LL_DFPQX4 \sa21_reg[6]  ( .D(N184), .CP(clk), .Q(sa21[6]) );
  HS65_LL_DFPQX4 \sa03_reg[5]  ( .D(N87), .CP(clk), .Q(sa03[5]) );
  HS65_LL_DFPQX4 \sa03_reg[6]  ( .D(N88), .CP(clk), .Q(sa03[6]) );
  HS65_LL_DFPQX4 \sa03_reg[7]  ( .D(N89), .CP(clk), .Q(sa03[7]) );
  HS65_LL_DFPQX4 \sa13_reg[6]  ( .D(N72), .CP(clk), .Q(sa13[6]) );
  HS65_LL_DFPQX4 \sa23_reg[6]  ( .D(N56), .CP(clk), .Q(sa23[6]) );
  HS65_LL_DFPQX4 \sa13_reg[7]  ( .D(N73), .CP(clk), .Q(sa13[7]) );
  HS65_LL_DFPQX4 \sa33_reg[6]  ( .D(N40), .CP(clk), .Q(sa33[6]) );
  HS65_LL_DFPQX4 \sa13_reg[3]  ( .D(N69), .CP(clk), .Q(sa13[3]) );
  HS65_LL_DFPQX4 \sa02_reg[6]  ( .D(N152), .CP(clk), .Q(sa02[6]) );
  HS65_LL_DFPQX4 \sa22_reg[5]  ( .D(N119), .CP(clk), .Q(sa22[5]) );
  HS65_LL_DFPQX4 \sa11_reg[3]  ( .D(N197), .CP(clk), .Q(sa11[3]) );
  HS65_LL_DFPQX4 \sa00_reg[0]  ( .D(N274), .CP(clk), .Q(sa00[0]) );
  HS65_LL_DFPQX4 \sa00_reg[3]  ( .D(N277), .CP(clk), .Q(sa00[3]) );
  HS65_LL_DFPQX4 \sa00_reg[1]  ( .D(N275), .CP(clk), .Q(sa00[1]) );
  HS65_LL_DFPQX4 \sa00_reg[4]  ( .D(N278), .CP(clk), .Q(sa00[4]) );
  HS65_LL_DFPQX4 \sa00_reg[5]  ( .D(N279), .CP(clk), .Q(sa00[5]) );
  HS65_LL_DFPQX4 \sa00_reg[6]  ( .D(N280), .CP(clk), .Q(sa00[6]) );
  HS65_LL_DFPQX4 \sa00_reg[7]  ( .D(N281), .CP(clk), .Q(sa00[7]) );
  HS65_LL_DFPQX4 \sa20_reg[7]  ( .D(N249), .CP(clk), .Q(sa20[7]) );
  HS65_LL_DFPQX4 \sa02_reg[5]  ( .D(N151), .CP(clk), .Q(sa02[5]) );
  HS65_LL_DFPQX4 \sa02_reg[7]  ( .D(N153), .CP(clk), .Q(sa02[7]) );
  HS65_LL_DFPQX4 \sa30_reg[6]  ( .D(N232), .CP(clk), .Q(sa30[6]) );
  HS65_LL_DFPQX4 \sa01_reg[1]  ( .D(N211), .CP(clk), .Q(sa01[1]) );
  HS65_LL_DFPQX4 \sa01_reg[2]  ( .D(N212), .CP(clk), .Q(sa01[2]) );
  HS65_LL_DFPQX4 \sa01_reg[4]  ( .D(N214), .CP(clk), .Q(sa01[4]) );
  HS65_LL_DFPQX4 \sa01_reg[3]  ( .D(N213), .CP(clk), .Q(sa01[3]) );
  HS65_LL_DFPQX4 \sa01_reg[5]  ( .D(N215), .CP(clk), .Q(sa01[5]) );
  HS65_LL_DFPQX4 \sa01_reg[6]  ( .D(N216), .CP(clk), .Q(sa01[6]) );
  HS65_LL_IVX18 U8573 ( .A(rst), .Z(N0) );
  HS65_LL_DFPQNX9 \dcnt_reg[3]  ( .D(n9113), .CP(clk), .QN(n2) );
  HS65_LLS_DFPQX18 \text_out_reg[16]  ( .D(N441), .CP(clk), .Q(text_out[16])
         );
  HS65_LLS_DFPQX18 \text_out_reg[15]  ( .D(N466), .CP(clk), .Q(text_out[15])
         );
  HS65_LLS_DFPQX18 \text_out_reg[105]  ( .D(N448), .CP(clk), .Q(text_out[105])
         );
  HS65_LLS_DFPQX18 \text_out_reg[4]  ( .D(N501), .CP(clk), .Q(text_out[4]) );
  HS65_LLS_DFPQX18 \text_out_reg[31]  ( .D(N402), .CP(clk), .Q(text_out[31])
         );
  HS65_LLS_DFPQX18 \text_out_reg[17]  ( .D(N440), .CP(clk), .Q(text_out[17])
         );
  HS65_LLS_DFPQX18 \text_out_reg[18]  ( .D(N439), .CP(clk), .Q(text_out[18])
         );
  HS65_LLS_DFPQX18 \text_out_reg[79]  ( .D(N450), .CP(clk), .Q(text_out[79])
         );
  HS65_LLS_DFPQX18 \text_out_reg[73]  ( .D(N456), .CP(clk), .Q(text_out[73])
         );
  HS65_LLS_DFPQX18 \text_out_reg[6]  ( .D(N499), .CP(clk), .Q(text_out[6]) );
  HS65_LLS_DFPQX18 \text_out_reg[23]  ( .D(N434), .CP(clk), .Q(text_out[23])
         );
  HS65_LLS_DFPQX18 \text_out_reg[56]  ( .D(N401), .CP(clk), .Q(text_out[56])
         );
  HS65_LLS_DFPQX18 \text_out_reg[0]  ( .D(N505), .CP(clk), .Q(text_out[0]) );
  HS65_LLS_DFPQX18 \text_out_reg[26]  ( .D(N407), .CP(clk), .Q(text_out[26])
         );
  HS65_LLS_DFPQX18 \text_out_reg[88]  ( .D(N393), .CP(clk), .Q(text_out[88])
         );
  HS65_LLS_DFPQX18 \text_out_reg[94]  ( .D(N387), .CP(clk), .Q(text_out[94])
         );
  HS65_LLS_DFPQX18 \text_out_reg[93]  ( .D(N388), .CP(clk), .Q(text_out[93])
         );
  HS65_LLS_DFPQX18 \text_out_reg[92]  ( .D(N389), .CP(clk), .Q(text_out[92])
         );
  HS65_LLS_DFPQX18 \text_out_reg[90]  ( .D(N391), .CP(clk), .Q(text_out[90])
         );
  HS65_LLS_DFPQX18 \text_out_reg[91]  ( .D(N390), .CP(clk), .Q(text_out[91])
         );
  HS65_LLS_DFPQX18 \text_out_reg[89]  ( .D(N392), .CP(clk), .Q(text_out[89])
         );
  HS65_LLS_DFPQX18 \text_out_reg[65]  ( .D(N488), .CP(clk), .Q(text_out[65])
         );
  HS65_LLS_DFPQX18 \text_out_reg[45]  ( .D(N460), .CP(clk), .Q(text_out[45])
         );
  HS65_LLS_DFPQX18 \text_out_reg[1]  ( .D(N504), .CP(clk), .Q(text_out[1]) );
  HS65_LLS_DFPQX18 \text_out_reg[43]  ( .D(N462), .CP(clk), .Q(text_out[43])
         );
  HS65_LLS_DFPQX18 \text_out_reg[82]  ( .D(N423), .CP(clk), .Q(text_out[82])
         );
  HS65_LLS_DFPQX18 \text_out_reg[60]  ( .D(N397), .CP(clk), .Q(text_out[60])
         );
  HS65_LLS_DFPQX18 \text_out_reg[59]  ( .D(N398), .CP(clk), .Q(text_out[59])
         );
  HS65_LLS_DFPQX18 \text_out_reg[62]  ( .D(N395), .CP(clk), .Q(text_out[62])
         );
  HS65_LLS_DFPQX18 \text_out_reg[52]  ( .D(N429), .CP(clk), .Q(text_out[52])
         );
  HS65_LLS_DFPQX18 \text_out_reg[46]  ( .D(N459), .CP(clk), .Q(text_out[46])
         );
  HS65_LLS_DFPQX18 \text_out_reg[121]  ( .D(N384), .CP(clk), .Q(text_out[121])
         );
  HS65_LLS_DFPQX18 \text_out_reg[126]  ( .D(N379), .CP(clk), .Q(text_out[126])
         );
  HS65_LLS_DFPQX18 \text_out_reg[125]  ( .D(N380), .CP(clk), .Q(text_out[125])
         );
  HS65_LLS_DFPQX18 \text_out_reg[124]  ( .D(N381), .CP(clk), .Q(text_out[124])
         );
  HS65_LLS_DFPQX18 \text_out_reg[123]  ( .D(N382), .CP(clk), .Q(text_out[123])
         );
  HS65_LLS_DFPQX18 \text_out_reg[120]  ( .D(N385), .CP(clk), .Q(text_out[120])
         );
  HS65_LLS_DFPQX18 \text_out_reg[122]  ( .D(N383), .CP(clk), .Q(text_out[122])
         );
  HS65_LLS_DFPQX18 \text_out_reg[21]  ( .D(N436), .CP(clk), .Q(text_out[21])
         );
  HS65_LLS_DFPQX18 \text_out_reg[118]  ( .D(N411), .CP(clk), .Q(text_out[118])
         );
  HS65_LLS_DFPQX18 \text_out_reg[75]  ( .D(N454), .CP(clk), .Q(text_out[75])
         );
  HS65_LLS_DFPQX18 \text_out_reg[55]  ( .D(N426), .CP(clk), .Q(text_out[55])
         );
  HS65_LLS_DFPQX18 \text_out_reg[110]  ( .D(N443), .CP(clk), .Q(text_out[110])
         );
  HS65_LLS_DFPQX18 \text_out_reg[109]  ( .D(N444), .CP(clk), .Q(text_out[109])
         );
  HS65_LLS_DFPQX18 \text_out_reg[53]  ( .D(N428), .CP(clk), .Q(text_out[53])
         );
  HS65_LLS_DFPQX18 \text_out_reg[10]  ( .D(N471), .CP(clk), .Q(text_out[10])
         );
  HS65_LLS_DFPQX18 \text_out_reg[12]  ( .D(N469), .CP(clk), .Q(text_out[12])
         );
  HS65_LLS_DFPQX18 \text_out_reg[97]  ( .D(N480), .CP(clk), .Q(text_out[97])
         );
  HS65_LLS_DFPQX18 \text_out_reg[25]  ( .D(N408), .CP(clk), .Q(text_out[25])
         );
  HS65_LLS_DFPQX18 \text_out_reg[27]  ( .D(N406), .CP(clk), .Q(text_out[27])
         );
  HS65_LLS_DFPQX18 \text_out_reg[30]  ( .D(N403), .CP(clk), .Q(text_out[30])
         );
  HS65_LLS_DFPQX18 \text_out_reg[29]  ( .D(N404), .CP(clk), .Q(text_out[29])
         );
  HS65_LLS_DFPQX18 \text_out_reg[14]  ( .D(N467), .CP(clk), .Q(text_out[14])
         );
  HS65_LLS_DFPQX18 \text_out_reg[13]  ( .D(N468), .CP(clk), .Q(text_out[13])
         );
  HS65_LLS_DFPQX18 \text_out_reg[77]  ( .D(N452), .CP(clk), .Q(text_out[77])
         );
  HS65_LLS_DFPQX18 \text_out_reg[78]  ( .D(N451), .CP(clk), .Q(text_out[78])
         );
  HS65_LLS_DFPQX18 \text_out_reg[22]  ( .D(N435), .CP(clk), .Q(text_out[22])
         );
  HS65_LLS_DFPQX18 \text_out_reg[19]  ( .D(N438), .CP(clk), .Q(text_out[19])
         );
  HS65_LLS_DFPQX18 \text_out_reg[127]  ( .D(N378), .CP(clk), .Q(text_out[127])
         );
  HS65_LLS_DFPQX18 \text_out_reg[113]  ( .D(N416), .CP(clk), .Q(text_out[113])
         );
  HS65_LLS_DFPQX18 \text_out_reg[86]  ( .D(N419), .CP(clk), .Q(text_out[86])
         );
  HS65_LLS_DFPQX18 \text_out_reg[54]  ( .D(N427), .CP(clk), .Q(text_out[54])
         );
  HS65_LLS_DFPQX18 \text_out_reg[20]  ( .D(N437), .CP(clk), .Q(text_out[20])
         );
  HS65_LLS_DFPQX18 \text_out_reg[107]  ( .D(N446), .CP(clk), .Q(text_out[107])
         );
  HS65_LLS_DFPQX18 \text_out_reg[63]  ( .D(N394), .CP(clk), .Q(text_out[63])
         );
  HS65_LLS_DFPQX18 \text_out_reg[51]  ( .D(N430), .CP(clk), .Q(text_out[51])
         );
  HS65_LLS_DFPQX18 \text_out_reg[9]  ( .D(N472), .CP(clk), .Q(text_out[9]) );
  HS65_LLS_DFPQX18 \text_out_reg[84]  ( .D(N421), .CP(clk), .Q(text_out[84])
         );
  HS65_LLS_DFPQX18 \text_out_reg[102]  ( .D(N475), .CP(clk), .Q(text_out[102])
         );
  HS65_LLS_DFPQX18 \text_out_reg[28]  ( .D(N405), .CP(clk), .Q(text_out[28])
         );
  HS65_LLS_DFPQX18 \text_out_reg[5]  ( .D(N500), .CP(clk), .Q(text_out[5]) );
  HS65_LLS_DFPQX18 \text_out_reg[44]  ( .D(N461), .CP(clk), .Q(text_out[44])
         );
  HS65_LLS_DFPQX18 \text_out_reg[116]  ( .D(N413), .CP(clk), .Q(text_out[116])
         );
  HS65_LLS_DFPQX18 \text_out_reg[85]  ( .D(N420), .CP(clk), .Q(text_out[85])
         );
  HS65_LLS_DFPQX18 \text_out_reg[101]  ( .D(N476), .CP(clk), .Q(text_out[101])
         );
  HS65_LLS_DFPQX18 \text_out_reg[48]  ( .D(N433), .CP(clk), .Q(text_out[48])
         );
  HS65_LLS_DFPQX18 \text_out_reg[119]  ( .D(N410), .CP(clk), .Q(text_out[119])
         );
  HS65_LLS_DFPQX18 \text_out_reg[76]  ( .D(N453), .CP(clk), .Q(text_out[76])
         );
  HS65_LLS_DFPQX18 \text_out_reg[61]  ( .D(N396), .CP(clk), .Q(text_out[61])
         );
  HS65_LLS_DFPQX18 \text_out_reg[58]  ( .D(N399), .CP(clk), .Q(text_out[58])
         );
  HS65_LLS_DFPQX18 \text_out_reg[57]  ( .D(N400), .CP(clk), .Q(text_out[57])
         );
  HS65_LLS_DFPQX18 \text_out_reg[49]  ( .D(N432), .CP(clk), .Q(text_out[49])
         );
  HS65_LLS_DFPQX18 \text_out_reg[11]  ( .D(N470), .CP(clk), .Q(text_out[11])
         );
  HS65_LLS_DFPQX18 \text_out_reg[117]  ( .D(N412), .CP(clk), .Q(text_out[117])
         );
  HS65_LLS_DFPQX18 \text_out_reg[83]  ( .D(N422), .CP(clk), .Q(text_out[83])
         );
  HS65_LLS_DFPQX18 \text_out_reg[40]  ( .D(N465), .CP(clk), .Q(text_out[40])
         );
  HS65_LLS_DFPQX18 \text_out_reg[96]  ( .D(N481), .CP(clk), .Q(text_out[96])
         );
  HS65_LLS_DFPQX18 \text_out_reg[24]  ( .D(N409), .CP(clk), .Q(text_out[24])
         );
  HS65_LLS_DFPQX18 \text_out_reg[108]  ( .D(N445), .CP(clk), .Q(text_out[108])
         );
  HS65_LLS_DFPQX18 \text_out_reg[47]  ( .D(N458), .CP(clk), .Q(text_out[47])
         );
  HS65_LLS_DFPQX18 \text_out_reg[106]  ( .D(N447), .CP(clk), .Q(text_out[106])
         );
  HS65_LLS_DFPQX18 \text_out_reg[37]  ( .D(N492), .CP(clk), .Q(text_out[37])
         );
  HS65_LLS_DFPQX18 \text_out_reg[69]  ( .D(N484), .CP(clk), .Q(text_out[69])
         );
  HS65_LLS_DFPQX18 \text_out_reg[114]  ( .D(N415), .CP(clk), .Q(text_out[114])
         );
  HS65_LLS_DFPQX18 \text_out_reg[81]  ( .D(N424), .CP(clk), .Q(text_out[81])
         );
  HS65_LLS_DFPQX18 \text_out_reg[41]  ( .D(N464), .CP(clk), .Q(text_out[41])
         );
  HS65_LLS_DFPQX18 \text_out_reg[98]  ( .D(N479), .CP(clk), .Q(text_out[98])
         );
  HS65_LLS_DFPQX18 \text_out_reg[3]  ( .D(N502), .CP(clk), .Q(text_out[3]) );
  HS65_LLS_DFPQX18 \text_out_reg[36]  ( .D(N493), .CP(clk), .Q(text_out[36])
         );
  HS65_LLS_DFPQX18 \text_out_reg[70]  ( .D(N483), .CP(clk), .Q(text_out[70])
         );
  HS65_LLS_DFPQX18 \text_out_reg[100]  ( .D(N477), .CP(clk), .Q(text_out[100])
         );
  HS65_LLS_DFPQX18 \text_out_reg[38]  ( .D(N491), .CP(clk), .Q(text_out[38])
         );
  HS65_LLS_DFPQX18 \text_out_reg[68]  ( .D(N485), .CP(clk), .Q(text_out[68])
         );
  HS65_LLS_DFPQX18 \text_out_reg[111]  ( .D(N442), .CP(clk), .Q(text_out[111])
         );
  HS65_LLS_DFPQX18 \text_out_reg[35]  ( .D(N494), .CP(clk), .Q(text_out[35])
         );
  HS65_LLS_DFPQX18 \text_out_reg[64]  ( .D(N489), .CP(clk), .Q(text_out[64])
         );
  HS65_LLS_DFPQX18 \text_out_reg[42]  ( .D(N463), .CP(clk), .Q(text_out[42])
         );
  HS65_LLS_DFPQX18 \text_out_reg[104]  ( .D(N449), .CP(clk), .Q(text_out[104])
         );
  HS65_LLS_DFPQX18 \text_out_reg[32]  ( .D(N497), .CP(clk), .Q(text_out[32])
         );
  HS65_LLS_DFPQX18 \text_out_reg[67]  ( .D(N486), .CP(clk), .Q(text_out[67])
         );
  HS65_LLS_DFPQX18 \text_out_reg[115]  ( .D(N414), .CP(clk), .Q(text_out[115])
         );
  HS65_LLS_DFPQX18 \text_out_reg[87]  ( .D(N418), .CP(clk), .Q(text_out[87])
         );
  HS65_LLS_DFPQX18 \text_out_reg[34]  ( .D(N495), .CP(clk), .Q(text_out[34])
         );
  HS65_LLS_DFPQX18 \text_out_reg[66]  ( .D(N487), .CP(clk), .Q(text_out[66])
         );
  HS65_LLS_DFPQX18 \text_out_reg[99]  ( .D(N478), .CP(clk), .Q(text_out[99])
         );
  HS65_LLS_DFPQX18 \text_out_reg[2]  ( .D(N503), .CP(clk), .Q(text_out[2]) );
  HS65_LLS_DFPQX18 \text_out_reg[39]  ( .D(N490), .CP(clk), .Q(text_out[39])
         );
  HS65_LLS_DFPQX18 \text_out_reg[74]  ( .D(N455), .CP(clk), .Q(text_out[74])
         );
  HS65_LLS_DFPQX18 \text_out_reg[72]  ( .D(N457), .CP(clk), .Q(text_out[72])
         );
  HS65_LLS_DFPQX18 \text_out_reg[112]  ( .D(N417), .CP(clk), .Q(text_out[112])
         );
  HS65_LLS_DFPQX18 \text_out_reg[80]  ( .D(N425), .CP(clk), .Q(text_out[80])
         );
  HS65_LLS_DFPQX18 \text_out_reg[50]  ( .D(N431), .CP(clk), .Q(text_out[50])
         );
  HS65_LLS_DFPQX18 \text_out_reg[8]  ( .D(N473), .CP(clk), .Q(text_out[8]) );
  HS65_LLS_DFPQX18 \text_out_reg[71]  ( .D(N482), .CP(clk), .Q(text_out[71])
         );
  HS65_LLS_DFPQX18 \text_out_reg[103]  ( .D(N474), .CP(clk), .Q(text_out[103])
         );
  HS65_LLS_DFPQX18 \text_out_reg[7]  ( .D(N498), .CP(clk), .Q(text_out[7]) );
  HS65_LLS_DFPQX18 \text_out_reg[33]  ( .D(N496), .CP(clk), .Q(text_out[33])
         );
  HS65_LLS_DFPQX18 \text_out_reg[95]  ( .D(N386), .CP(clk), .Q(text_out[95])
         );
  HS65_LLS_DFPQX18 done_reg ( .D(N23), .CP(clk), .Q(done) );
  HS65_LL_DFPHQX4 \text_in_r_reg[126]  ( .D(text_in[126]), .E(n9116), .CP(clk), 
        .Q(text_in_r[126]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[125]  ( .D(text_in[125]), .E(n9115), .CP(clk), 
        .Q(text_in_r[125]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[124]  ( .D(text_in[124]), .E(n9120), .CP(clk), 
        .Q(text_in_r[124]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[123]  ( .D(text_in[123]), .E(n9116), .CP(clk), 
        .Q(text_in_r[123]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[122]  ( .D(text_in[122]), .E(n9119), .CP(clk), 
        .Q(text_in_r[122]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[121]  ( .D(text_in[121]), .E(ld), .CP(clk), 
        .Q(text_in_r[121]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[120]  ( .D(text_in[120]), .E(n9116), .CP(clk), 
        .Q(text_in_r[120]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[119]  ( .D(text_in[119]), .E(n9115), .CP(clk), 
        .Q(text_in_r[119]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[118]  ( .D(text_in[118]), .E(n9120), .CP(clk), 
        .Q(text_in_r[118]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[117]  ( .D(text_in[117]), .E(n9116), .CP(clk), 
        .Q(text_in_r[117]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[116]  ( .D(text_in[116]), .E(n9119), .CP(clk), 
        .Q(text_in_r[116]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[115]  ( .D(text_in[115]), .E(ld), .CP(clk), 
        .Q(text_in_r[115]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[114]  ( .D(text_in[114]), .E(n9116), .CP(clk), 
        .Q(text_in_r[114]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[113]  ( .D(text_in[113]), .E(n9120), .CP(clk), 
        .Q(text_in_r[113]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[112]  ( .D(text_in[112]), .E(ld), .CP(clk), 
        .Q(text_in_r[112]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[111]  ( .D(text_in[111]), .E(n9116), .CP(clk), 
        .Q(text_in_r[111]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[110]  ( .D(text_in[110]), .E(n9115), .CP(clk), 
        .Q(text_in_r[110]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[109]  ( .D(text_in[109]), .E(n9150), .CP(clk), 
        .Q(text_in_r[109]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[108]  ( .D(text_in[108]), .E(n9116), .CP(clk), 
        .Q(text_in_r[108]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[107]  ( .D(text_in[107]), .E(n9119), .CP(clk), 
        .Q(text_in_r[107]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[106]  ( .D(text_in[106]), .E(n9120), .CP(clk), 
        .Q(text_in_r[106]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[105]  ( .D(text_in[105]), .E(n9116), .CP(clk), 
        .Q(text_in_r[105]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[104]  ( .D(text_in[104]), .E(n9115), .CP(clk), 
        .Q(text_in_r[104]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[103]  ( .D(text_in[103]), .E(n9150), .CP(clk), 
        .Q(text_in_r[103]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[102]  ( .D(text_in[102]), .E(n9116), .CP(clk), 
        .Q(text_in_r[102]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[101]  ( .D(text_in[101]), .E(n9119), .CP(clk), 
        .Q(text_in_r[101]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[100]  ( .D(text_in[100]), .E(n9150), .CP(clk), 
        .Q(text_in_r[100]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[99]  ( .D(text_in[99]), .E(n9116), .CP(clk), 
        .Q(text_in_r[99]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[98]  ( .D(text_in[98]), .E(n9115), .CP(clk), 
        .Q(text_in_r[98]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[97]  ( .D(text_in[97]), .E(n9150), .CP(clk), 
        .Q(text_in_r[97]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[96]  ( .D(text_in[96]), .E(n9116), .CP(clk), 
        .Q(text_in_r[96]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[95]  ( .D(text_in[95]), .E(n9119), .CP(clk), 
        .Q(text_in_r[95]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[94]  ( .D(text_in[94]), .E(n9150), .CP(clk), 
        .Q(text_in_r[94]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[93]  ( .D(text_in[93]), .E(n9116), .CP(clk), 
        .Q(text_in_r[93]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[92]  ( .D(text_in[92]), .E(n9120), .CP(clk), 
        .Q(text_in_r[92]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[91]  ( .D(text_in[91]), .E(n9150), .CP(clk), 
        .Q(text_in_r[91]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[90]  ( .D(text_in[90]), .E(n9116), .CP(clk), 
        .Q(text_in_r[90]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[89]  ( .D(text_in[89]), .E(n9115), .CP(clk), 
        .Q(text_in_r[89]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[88]  ( .D(text_in[88]), .E(n9150), .CP(clk), 
        .Q(text_in_r[88]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[87]  ( .D(text_in[87]), .E(n9116), .CP(clk), 
        .Q(text_in_r[87]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[86]  ( .D(text_in[86]), .E(n9119), .CP(clk), 
        .Q(text_in_r[86]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[85]  ( .D(text_in[85]), .E(n9150), .CP(clk), 
        .Q(text_in_r[85]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[84]  ( .D(text_in[84]), .E(n9116), .CP(clk), 
        .Q(text_in_r[84]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[83]  ( .D(text_in[83]), .E(n9115), .CP(clk), 
        .Q(text_in_r[83]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[82]  ( .D(text_in[82]), .E(n9150), .CP(clk), 
        .Q(text_in_r[82]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[81]  ( .D(text_in[81]), .E(n9116), .CP(clk), 
        .Q(text_in_r[81]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[80]  ( .D(text_in[80]), .E(n9119), .CP(clk), 
        .Q(text_in_r[80]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[79]  ( .D(text_in[79]), .E(n9150), .CP(clk), 
        .Q(text_in_r[79]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[78]  ( .D(text_in[78]), .E(n9116), .CP(clk), 
        .Q(text_in_r[78]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[77]  ( .D(text_in[77]), .E(n9115), .CP(clk), 
        .Q(text_in_r[77]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[76]  ( .D(text_in[76]), .E(n9150), .CP(clk), 
        .Q(text_in_r[76]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[75]  ( .D(text_in[75]), .E(n9116), .CP(clk), 
        .Q(text_in_r[75]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[74]  ( .D(text_in[74]), .E(n9119), .CP(clk), 
        .Q(text_in_r[74]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[73]  ( .D(text_in[73]), .E(n9150), .CP(clk), 
        .Q(text_in_r[73]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[72]  ( .D(text_in[72]), .E(n9116), .CP(clk), 
        .Q(text_in_r[72]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[71]  ( .D(text_in[71]), .E(n9120), .CP(clk), 
        .Q(text_in_r[71]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[70]  ( .D(text_in[70]), .E(n9150), .CP(clk), 
        .Q(text_in_r[70]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[69]  ( .D(text_in[69]), .E(n9117), .CP(clk), 
        .Q(text_in_r[69]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[68]  ( .D(text_in[68]), .E(n9115), .CP(clk), 
        .Q(text_in_r[68]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[67]  ( .D(text_in[67]), .E(n9150), .CP(clk), 
        .Q(text_in_r[67]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[66]  ( .D(text_in[66]), .E(n9117), .CP(clk), 
        .Q(text_in_r[66]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[65]  ( .D(text_in[65]), .E(n9119), .CP(clk), 
        .Q(text_in_r[65]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[64]  ( .D(text_in[64]), .E(n9115), .CP(clk), 
        .Q(text_in_r[64]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[63]  ( .D(text_in[63]), .E(n9150), .CP(clk), 
        .Q(text_in_r[63]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[62]  ( .D(text_in[62]), .E(n9117), .CP(clk), 
        .Q(text_in_r[62]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[61]  ( .D(text_in[61]), .E(n9121), .CP(clk), 
        .Q(text_in_r[61]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[60]  ( .D(text_in[60]), .E(n9117), .CP(clk), 
        .Q(text_in_r[60]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[59]  ( .D(text_in[59]), .E(n9119), .CP(clk), 
        .Q(text_in_r[59]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[58]  ( .D(text_in[58]), .E(n9121), .CP(clk), 
        .Q(text_in_r[58]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[57]  ( .D(text_in[57]), .E(n9117), .CP(clk), 
        .Q(text_in_r[57]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[56]  ( .D(text_in[56]), .E(n9115), .CP(clk), 
        .Q(text_in_r[56]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[55]  ( .D(text_in[55]), .E(n9119), .CP(clk), 
        .Q(text_in_r[55]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[54]  ( .D(text_in[54]), .E(n9121), .CP(clk), 
        .Q(text_in_r[54]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[53]  ( .D(text_in[53]), .E(n9117), .CP(clk), 
        .Q(text_in_r[53]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[52]  ( .D(text_in[52]), .E(n9121), .CP(clk), 
        .Q(text_in_r[52]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[51]  ( .D(text_in[51]), .E(n9117), .CP(clk), 
        .Q(text_in_r[51]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[50]  ( .D(text_in[50]), .E(n9120), .CP(clk), 
        .Q(text_in_r[50]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[49]  ( .D(text_in[49]), .E(n9119), .CP(clk), 
        .Q(text_in_r[49]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[48]  ( .D(text_in[48]), .E(n9115), .CP(clk), 
        .Q(text_in_r[48]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[47]  ( .D(text_in[47]), .E(n9119), .CP(clk), 
        .Q(text_in_r[47]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[46]  ( .D(text_in[46]), .E(n9115), .CP(clk), 
        .Q(text_in_r[46]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[45]  ( .D(text_in[45]), .E(n9119), .CP(clk), 
        .Q(text_in_r[45]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[44]  ( .D(text_in[44]), .E(n9120), .CP(clk), 
        .Q(text_in_r[44]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[43]  ( .D(text_in[43]), .E(n9115), .CP(clk), 
        .Q(text_in_r[43]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[42]  ( .D(text_in[42]), .E(n9119), .CP(clk), 
        .Q(text_in_r[42]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[41]  ( .D(text_in[41]), .E(n9120), .CP(clk), 
        .Q(text_in_r[41]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[40]  ( .D(text_in[40]), .E(n9120), .CP(clk), 
        .Q(text_in_r[40]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[30]  ( .D(text_in[30]), .E(n9120), .CP(clk), 
        .Q(text_in_r[30]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[127]  ( .D(text_in[127]), .E(n9150), .CP(clk), 
        .Q(text_in_r[127]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[39]  ( .D(text_in[39]), .E(n9121), .CP(clk), 
        .Q(text_in_r[39]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[38]  ( .D(text_in[38]), .E(n9117), .CP(clk), 
        .Q(text_in_r[38]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[37]  ( .D(text_in[37]), .E(n9115), .CP(clk), 
        .Q(text_in_r[37]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[36]  ( .D(text_in[36]), .E(n9119), .CP(clk), 
        .Q(text_in_r[36]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[35]  ( .D(text_in[35]), .E(n9121), .CP(clk), 
        .Q(text_in_r[35]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[34]  ( .D(text_in[34]), .E(n9117), .CP(clk), 
        .Q(text_in_r[34]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[33]  ( .D(text_in[33]), .E(n9121), .CP(clk), 
        .Q(text_in_r[33]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[32]  ( .D(text_in[32]), .E(n9117), .CP(clk), 
        .Q(text_in_r[32]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[31]  ( .D(text_in[31]), .E(n9115), .CP(clk), 
        .Q(text_in_r[31]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[29]  ( .D(text_in[29]), .E(n9119), .CP(clk), 
        .Q(text_in_r[29]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[28]  ( .D(text_in[28]), .E(n9121), .CP(clk), 
        .Q(text_in_r[28]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[27]  ( .D(text_in[27]), .E(n9117), .CP(clk), 
        .Q(text_in_r[27]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[26]  ( .D(text_in[26]), .E(n9120), .CP(clk), 
        .Q(text_in_r[26]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[25]  ( .D(text_in[25]), .E(n9121), .CP(clk), 
        .Q(text_in_r[25]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[24]  ( .D(text_in[24]), .E(n9117), .CP(clk), 
        .Q(text_in_r[24]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[23]  ( .D(text_in[23]), .E(n9115), .CP(clk), 
        .Q(text_in_r[23]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[22]  ( .D(text_in[22]), .E(n9121), .CP(clk), 
        .Q(text_in_r[22]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[21]  ( .D(text_in[21]), .E(n9117), .CP(clk), 
        .Q(text_in_r[21]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[20]  ( .D(text_in[20]), .E(n9121), .CP(clk), 
        .Q(text_in_r[20]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[19]  ( .D(text_in[19]), .E(n9117), .CP(clk), 
        .Q(text_in_r[19]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[18]  ( .D(text_in[18]), .E(n9119), .CP(clk), 
        .Q(text_in_r[18]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[17]  ( .D(text_in[17]), .E(n9115), .CP(clk), 
        .Q(text_in_r[17]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[16]  ( .D(text_in[16]), .E(n9121), .CP(clk), 
        .Q(text_in_r[16]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[15]  ( .D(text_in[15]), .E(n9117), .CP(clk), 
        .Q(text_in_r[15]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[14]  ( .D(text_in[14]), .E(n9119), .CP(clk), 
        .Q(text_in_r[14]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[13]  ( .D(text_in[13]), .E(n9121), .CP(clk), 
        .Q(text_in_r[13]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[12]  ( .D(text_in[12]), .E(n9117), .CP(clk), 
        .Q(text_in_r[12]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[11]  ( .D(text_in[11]), .E(n9115), .CP(clk), 
        .Q(text_in_r[11]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[10]  ( .D(text_in[10]), .E(n9121), .CP(clk), 
        .Q(text_in_r[10]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[9]  ( .D(text_in[9]), .E(n9117), .CP(clk), 
        .Q(text_in_r[9]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[8]  ( .D(text_in[8]), .E(n9119), .CP(clk), 
        .Q(text_in_r[8]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[7]  ( .D(text_in[7]), .E(n9121), .CP(clk), 
        .Q(text_in_r[7]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[6]  ( .D(text_in[6]), .E(n9117), .CP(clk), 
        .Q(text_in_r[6]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[5]  ( .D(text_in[5]), .E(n9120), .CP(clk), 
        .Q(text_in_r[5]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[4]  ( .D(text_in[4]), .E(n9121), .CP(clk), 
        .Q(text_in_r[4]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[3]  ( .D(text_in[3]), .E(n9117), .CP(clk), 
        .Q(text_in_r[3]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[2]  ( .D(text_in[2]), .E(n9115), .CP(clk), 
        .Q(text_in_r[2]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[1]  ( .D(text_in[1]), .E(n9121), .CP(clk), 
        .Q(text_in_r[1]) );
  HS65_LL_DFPHQX4 \text_in_r_reg[0]  ( .D(text_in[0]), .E(n9117), .CP(clk), 
        .Q(text_in_r[0]) );
  HS65_LL_DFPQNX9 ld_r_reg ( .D(n9121), .CP(clk), .QN(n9136) );
  HS65_LL_IVX7 U9537 ( .A(n9118), .Z(n9115) );
  HS65_LL_IVX9 U9538 ( .A(n9143), .Z(n9116) );
  HS65_LL_IVX9 U9539 ( .A(n9143), .Z(n9117) );
  HS65_LL_IVX2 U9540 ( .A(ld), .Z(n9118) );
  HS65_LL_IVX7 U9541 ( .A(n9118), .Z(n9119) );
  HS65_LL_IVX2 U9542 ( .A(n9118), .Z(n9120) );
  HS65_LL_IVX9 U9543 ( .A(n9118), .Z(n9121) );
  HS65_LL_AND2X4 U9544 ( .A(n5741), .B(n5740), .Z(n4481) );
  HS65_LL_AND2X4 U9545 ( .A(n7333), .B(n7332), .Z(n6074) );
  HS65_LL_AND2X4 U9546 ( .A(n5803), .B(n5802), .Z(n4521) );
  HS65_LL_AND2X4 U9547 ( .A(n7395), .B(n7394), .Z(n6114) );
  HS65_LL_AND2X4 U9548 ( .A(n5877), .B(n5863), .Z(n4589) );
  HS65_LL_AND2X4 U9549 ( .A(n7528), .B(n7514), .Z(n6199) );
  HS65_LL_AND2X4 U9550 ( .A(n7460), .B(n7457), .Z(n6182) );
  HS65_LL_AND2X4 U9551 ( .A(n5936), .B(n5922), .Z(n4606) );
  HS65_LL_AND2X4 U9552 ( .A(n9049), .B(n9034), .Z(n7699) );
  HS65_LL_AND2X4 U9553 ( .A(n9107), .B(n9092), .Z(n7737) );
  HS65_LL_IVX9 U9554 ( .A(n7550), .Z(n94) );
  HS65_LLS_XNOR2X6 U9555 ( .A(n2817), .B(n2793), .Z(n4364) );
  HS65_LLS_XNOR2X6 U9556 ( .A(n315), .B(n2750), .Z(n2619) );
  HS65_LLS_XNOR2X6 U9557 ( .A(n2809), .B(n2785), .Z(n5957) );
  HS65_LLS_XNOR2X6 U9558 ( .A(n2703), .B(n2653), .Z(n2660) );
  HS65_LLS_XNOR2X6 U9559 ( .A(n2652), .B(n2733), .Z(n2702) );
  HS65_LLS_XOR2X6 U9560 ( .A(n2718), .B(n2672), .Z(n2677) );
  HS65_LLS_XOR2X6 U9561 ( .A(n2674), .B(n183), .Z(n2716) );
  HS65_LLS_XOR2X6 U9562 ( .A(n2801), .B(n573), .Z(n7550) );
  HS65_LLS_XNOR2X6 U9563 ( .A(n2653), .B(n2654), .Z(n2648) );
  HS65_LLS_XOR2X6 U9564 ( .A(n2703), .B(n2628), .Z(n2731) );
  HS65_LLS_XOR2X6 U9565 ( .A(n2718), .B(n2628), .Z(n2744) );
  HS65_LLS_XNOR2X6 U9566 ( .A(n2817), .B(n4347), .Z(n4427) );
  HS65_LLS_XNOR2X6 U9567 ( .A(n2809), .B(n5940), .Z(n6020) );
  HS65_LLS_XOR2X6 U9568 ( .A(n2801), .B(n7532), .Z(n7609) );
  HS65_LL_IVX9 U9569 ( .A(n4347), .Z(n7) );
  HS65_LL_IVX9 U9570 ( .A(n5940), .Z(n52) );
  HS65_LLS_XOR2X6 U9571 ( .A(n3001), .B(n7546), .Z(n7543) );
  HS65_LLS_XOR2X6 U9572 ( .A(n2672), .B(n2654), .Z(n2671) );
  HS65_LLS_XNOR2X6 U9573 ( .A(n3009), .B(n272), .Z(n5951) );
  HS65_LLS_XNOR2X6 U9574 ( .A(n3212), .B(n447), .Z(n4358) );
  HS65_LL_IVX9 U9575 ( .A(n5968), .Z(n272) );
  HS65_LL_IVX9 U9576 ( .A(n4375), .Z(n447) );
  HS65_LL_IVX9 U9577 ( .A(n2745), .Z(n183) );
  HS65_LL_NOR4ABX2 U9578 ( .A(n8325), .B(n7944), .C(n8315), .D(n8042), .Z(
        n8496) );
  HS65_LL_NOR4ABX2 U9579 ( .A(n2847), .B(n3958), .C(n3968), .D(n4025), .Z(
        n4287) );
  HS65_LL_NOR4ABX2 U9580 ( .A(n2877), .B(n3938), .C(n3948), .D(n4002), .Z(
        n4228) );
  HS65_LL_NOR4ABX2 U9581 ( .A(n2907), .B(n3019), .C(n3227), .D(n3237), .Z(
        n3539) );
  HS65_LL_NOR4ABX2 U9582 ( .A(n2987), .B(n3170), .C(n3356), .D(n3366), .Z(
        n3773) );
  HS65_LL_NOR4ABX2 U9583 ( .A(n2259), .B(n2517), .C(n2508), .D(n2530), .Z(
        n2552) );
  HS65_LL_NOR4ABX2 U9584 ( .A(n1883), .B(n2141), .C(n2132), .D(n2154), .Z(
        n2176) );
  HS65_LL_NOR4ABX2 U9585 ( .A(n1507), .B(n1765), .C(n1756), .D(n1778), .Z(
        n1800) );
  HS65_LL_NOR4ABX2 U9586 ( .A(n1131), .B(n1389), .C(n1380), .D(n1402), .Z(
        n1424) );
  HS65_LL_NOR4ABX2 U9587 ( .A(n97), .B(n8428), .C(n8439), .D(n8015), .Z(n8754)
         );
  HS65_LL_IVX9 U9588 ( .A(n8162), .Z(n97) );
  HS65_LL_NOR3AX2 U9589 ( .A(n6264), .B(n6289), .C(n6135), .Z(n6600) );
  HS65_LL_NOR3AX2 U9590 ( .A(n4671), .B(n4696), .C(n4542), .Z(n5007) );
  HS65_LL_NOR3AX2 U9591 ( .A(n8375), .B(n8386), .C(n8138), .Z(n8672) );
  HS65_LL_NOR3AX2 U9592 ( .A(n8427), .B(n8438), .C(n8161), .Z(n8762) );
  HS65_LL_NAND2X7 U9593 ( .A(n913), .B(n896), .Z(n2332) );
  HS65_LL_NAND2X7 U9594 ( .A(n872), .B(n855), .Z(n1204) );
  HS65_LL_NAND2X7 U9595 ( .A(n831), .B(n814), .Z(n1580) );
  HS65_LL_NAND2X7 U9596 ( .A(n790), .B(n773), .Z(n1956) );
  HS65_LL_NOR4ABX2 U9597 ( .A(n3892), .B(n4050), .C(n4051), .D(n3920), .Z(
        n4044) );
  HS65_LL_NOR4ABX2 U9598 ( .A(n2864), .B(n2943), .C(n3071), .D(n3081), .Z(
        n3413) );
  HS65_LL_IVX9 U9599 ( .A(n2777), .Z(n573) );
  HS65_LL_NOR4ABX2 U9600 ( .A(n577), .B(n8376), .C(n8387), .D(n8002), .Z(n8662) );
  HS65_LL_IVX9 U9601 ( .A(n8139), .Z(n577) );
  HS65_LL_NOR3AX2 U9602 ( .A(n8314), .B(n8326), .C(n8041), .Z(n8530) );
  HS65_LL_NOR3AX2 U9603 ( .A(n3226), .B(n3238), .C(n3018), .Z(n3589) );
  HS65_LL_NOR3AX2 U9604 ( .A(n8068), .B(n8092), .C(n7973), .Z(n8228) );
  HS65_LL_NOR3AX2 U9605 ( .A(n3301), .B(n3313), .C(n3143), .Z(n3706) );
  HS65_LL_IVX9 U9606 ( .A(n2898), .Z(n315) );
  HS65_LL_IVX9 U9607 ( .A(n2056), .Z(n764) );
  HS65_LL_IVX9 U9608 ( .A(n2432), .Z(n887) );
  HS65_LL_IVX9 U9609 ( .A(n1304), .Z(n846) );
  HS65_LL_IVX9 U9610 ( .A(n1680), .Z(n805) );
  HS65_LL_IVX9 U9611 ( .A(n3717), .Z(n657) );
  HS65_LL_IVX9 U9612 ( .A(n8240), .Z(n388) );
  HS65_LL_IVX9 U9613 ( .A(n2733), .Z(n184) );
  HS65_LLS_XNOR2X6 U9614 ( .A(n3001), .B(n2753), .Z(n7582) );
  HS65_LL_IVX9 U9615 ( .A(n8629), .Z(n346) );
  HS65_LL_IVX9 U9616 ( .A(n3935), .Z(n647) );
  HS65_LL_IVX9 U9617 ( .A(n3973), .Z(n434) );
  HS65_LLS_XOR2X6 U9618 ( .A(n3009), .B(n2761), .Z(n5992) );
  HS65_LLS_XOR2X6 U9619 ( .A(n3212), .B(n2769), .Z(n4399) );
  HS65_LL_NOR4ABX2 U9620 ( .A(n4080), .B(n4081), .C(n3907), .D(n3987), .Z(
        n4076) );
  HS65_LL_NOR3AX2 U9621 ( .A(n3019), .B(n3020), .C(n2909), .Z(n3015) );
  HS65_LL_IVX9 U9622 ( .A(n9144), .Z(n9138) );
  HS65_LL_IVX9 U9623 ( .A(n9144), .Z(n9139) );
  HS65_LL_IVX9 U9624 ( .A(n9144), .Z(n9137) );
  HS65_LL_IVX9 U9625 ( .A(n5012), .Z(n38) );
  HS65_LL_IVX9 U9626 ( .A(n6605), .Z(n560) );
  HS65_LL_IVX9 U9627 ( .A(n3477), .Z(n208) );
  HS65_LL_IVX9 U9628 ( .A(n3832), .Z(n426) );
  HS65_LL_IVX9 U9629 ( .A(n3601), .Z(n171) );
  HS65_LL_IVX9 U9630 ( .A(n6959), .Z(n308) );
  HS65_LL_IVX9 U9631 ( .A(n6844), .Z(n80) );
  HS65_LL_IVX9 U9632 ( .A(n5252), .Z(n266) );
  HS65_LL_IVX9 U9633 ( .A(n5367), .Z(n483) );
  HS65_LL_IVX9 U9634 ( .A(n6726), .Z(n517) );
  HS65_LL_IVX9 U9635 ( .A(n5134), .Z(n693) );
  HS65_LL_IVX9 U9636 ( .A(n8542), .Z(n339) );
  HS65_LL_IVX9 U9637 ( .A(n8677), .Z(n608) );
  HS65_LL_IVX9 U9638 ( .A(n8767), .Z(n128) );
  HS65_LL_IVX9 U9639 ( .A(n9143), .Z(n9141) );
  HS65_LL_IVX9 U9640 ( .A(n9143), .Z(n9140) );
  HS65_LL_IVX9 U9641 ( .A(n9143), .Z(n9142) );
  HS65_LL_NAND3X5 U9642 ( .A(n8758), .B(n8759), .C(n7909), .Z(n8757) );
  HS65_LL_NAND3X5 U9643 ( .A(n8668), .B(n8669), .C(n7811), .Z(n8667) );
  HS65_LL_NAND3X5 U9644 ( .A(n8197), .B(n8198), .C(n8199), .Z(n8196) );
  HS65_LL_NAND3X5 U9645 ( .A(n6834), .B(n6835), .C(n6836), .Z(n6833) );
  HS65_LL_NAND3X5 U9646 ( .A(n5242), .B(n5243), .C(n5244), .Z(n5241) );
  HS65_LL_NAND3X5 U9647 ( .A(n5357), .B(n5358), .C(n5359), .Z(n5356) );
  HS65_LL_NAND3X5 U9648 ( .A(n5124), .B(n5125), .C(n5126), .Z(n5123) );
  HS65_LL_NAND3X5 U9649 ( .A(n6949), .B(n6950), .C(n6951), .Z(n6948) );
  HS65_LL_NAND3X5 U9650 ( .A(n6716), .B(n6717), .C(n6718), .Z(n6715) );
  HS65_LL_IVX9 U9651 ( .A(n9135), .Z(n9124) );
  HS65_LL_IVX9 U9652 ( .A(n9136), .Z(n9123) );
  HS65_LL_IVX9 U9653 ( .A(n9134), .Z(n9126) );
  HS65_LL_IVX9 U9654 ( .A(n9136), .Z(n9122) );
  HS65_LL_IVX9 U9655 ( .A(n9135), .Z(n9125) );
  HS65_LL_IVX9 U9656 ( .A(n7086), .Z(n507) );
  HS65_LL_IVX9 U9657 ( .A(n5494), .Z(n683) );
  HS65_LL_IVX9 U9658 ( .A(n5537), .Z(n254) );
  HS65_LL_IVX9 U9659 ( .A(n5559), .Z(n471) );
  HS65_LL_IVX9 U9660 ( .A(n7151), .Z(n296) );
  HS65_LL_IVX9 U9661 ( .A(n7129), .Z(n72) );
  HS65_LL_IVX9 U9662 ( .A(n8481), .Z(n385) );
  HS65_LL_IVX9 U9663 ( .A(n7062), .Z(n550) );
  HS65_LL_IVX9 U9664 ( .A(n5470), .Z(n28) );
  HS65_LL_IVX9 U9665 ( .A(n8719), .Z(n598) );
  HS65_LL_IVX9 U9666 ( .A(n8809), .Z(n118) );
  HS65_LL_IVX9 U9667 ( .A(n3890), .Z(n217) );
  HS65_LLS_XNOR2X6 U9668 ( .A(n2722), .B(n2749), .Z(n2628) );
  HS65_LLS_XOR2X6 U9669 ( .A(n2757), .B(n2781), .Z(n7532) );
  HS65_LLS_XOR2X6 U9670 ( .A(n3005), .B(n2805), .Z(n7546) );
  HS65_LLS_XOR2X6 U9671 ( .A(n2630), .B(n2682), .Z(n2654) );
  HS65_LLS_XNOR2X6 U9672 ( .A(n2805), .B(n2781), .Z(n7576) );
  HS65_LLS_XNOR2X6 U9673 ( .A(n2797), .B(n2773), .Z(n4347) );
  HS65_LLS_XNOR2X6 U9674 ( .A(n2789), .B(n2765), .Z(n5940) );
  HS65_LLS_XNOR2X6 U9675 ( .A(n3207), .B(n2764), .Z(n5978) );
  HS65_LLS_XNOR2X6 U9676 ( .A(n3532), .B(n2772), .Z(n4385) );
  HS65_LLS_XNOR2X6 U9677 ( .A(n3004), .B(n2756), .Z(n7568) );
  HS65_LLS_XNOR2X6 U9678 ( .A(n2698), .B(n2641), .Z(n2649) );
  HS65_LLS_XNOR2X6 U9679 ( .A(n2818), .B(n2794), .Z(n4359) );
  HS65_LLS_XNOR2X6 U9680 ( .A(n3006), .B(n2758), .Z(n6003) );
  HS65_LLS_XNOR2X6 U9681 ( .A(n2806), .B(n2782), .Z(n5971) );
  HS65_LLS_XNOR2X6 U9682 ( .A(n2810), .B(n2786), .Z(n5952) );
  HS65_LLS_XNOR2X6 U9683 ( .A(n2751), .B(n2620), .Z(n7590) );
  HS65_LLS_XOR2X6 U9684 ( .A(n2630), .B(n404), .Z(n2695) );
  HS65_LL_NOR4ABX2 U9685 ( .A(n7739), .B(n7740), .C(n7741), .D(n7742), .Z(
        n2750) );
  HS65_LL_MX41X7 U9686 ( .D0(n362), .S0(n400), .D1(n394), .S1(n366), .D2(n367), 
        .S2(n387), .D3(n373), .S3(n393), .Z(n7741) );
  HS65_LL_MX41X7 U9687 ( .D0(n399), .S0(n368), .D1(n377), .S1(n383), .D2(n375), 
        .S2(n397), .D3(n370), .S3(n7743), .Z(n7742) );
  HS65_LL_NOR4ABX2 U9688 ( .A(n7744), .B(n7745), .C(n7746), .D(n7747), .Z(
        n7740) );
  HS65_LLS_XOR2X6 U9689 ( .A(n2757), .B(n316), .Z(n2616) );
  HS65_LLS_XNOR2X6 U9690 ( .A(n2820), .B(n231), .Z(n4351) );
  HS65_LLS_XNOR2X6 U9691 ( .A(n2812), .B(n53), .Z(n5944) );
  HS65_LL_NOR4ABX2 U9692 ( .A(n3656), .B(n3657), .C(n3658), .D(n3659), .Z(
        n2653) );
  HS65_LL_MX41X7 U9693 ( .D0(n661), .S0(n631), .D1(n630), .S1(n651), .D2(n652), 
        .S2(n628), .D3(n629), .S3(n3163), .Z(n3659) );
  HS65_LL_MX41X7 U9694 ( .D0(n633), .S0(n644), .D1(n627), .S1(n648), .D2(n624), 
        .S2(n645), .D3(n650), .S3(n625), .Z(n3658) );
  HS65_LL_AOI212X4 U9695 ( .A(n660), .B(n3660), .C(n626), .D(n3330), .E(n3661), 
        .Z(n3657) );
  HS65_LL_NOR4ABX2 U9696 ( .A(n8191), .B(n8192), .C(n8193), .D(n8194), .Z(
        n2753) );
  HS65_LL_MX41X7 U9697 ( .D0(n367), .S0(n387), .D1(n374), .S1(n386), .D2(n373), 
        .S2(n383), .D3(n393), .S3(n372), .Z(n8193) );
  HS65_LL_MX41X7 U9698 ( .D0(n392), .S0(n378), .D1(n376), .S1(n396), .D2(n395), 
        .S2(n377), .D3(n375), .S3(n7743), .Z(n8194) );
  HS65_LL_AOI212X4 U9699 ( .A(n391), .B(n8195), .C(n371), .D(n8110), .E(n8196), 
        .Z(n8192) );
  HS65_LLS_XOR2X6 U9700 ( .A(n3533), .B(n448), .Z(n4375) );
  HS65_LLS_XOR2X6 U9701 ( .A(n3208), .B(n273), .Z(n5968) );
  HS65_LLS_XOR2X6 U9702 ( .A(n2722), .B(n2682), .Z(n3218) );
  HS65_LL_NOR4ABX2 U9703 ( .A(n6828), .B(n6829), .C(n6830), .D(n6831), .Z(
        n2785) );
  HS65_LL_MX41X7 U9704 ( .D0(n63), .S0(n78), .D1(n77), .S1(n66), .D2(n73), 
        .S2(n65), .D3(n64), .S3(n6338), .Z(n6831) );
  HS65_LL_MX41X7 U9705 ( .D0(n57), .S0(n91), .D1(n90), .S1(n62), .D2(n89), 
        .S2(n59), .D3(n60), .S3(n76), .Z(n6830) );
  HS65_LL_AOI212X4 U9706 ( .A(n79), .B(n6832), .C(n58), .D(n6520), .E(n6833), 
        .Z(n6829) );
  HS65_LL_NOR4ABX2 U9707 ( .A(n5236), .B(n5237), .C(n5238), .D(n5239), .Z(
        n2793) );
  HS65_LL_MX41X7 U9708 ( .D0(n234), .S0(n264), .D1(n259), .S1(n235), .D2(n258), 
        .S2(n232), .D3(n233), .S3(n4757), .Z(n5239) );
  HS65_LL_MX41X7 U9709 ( .D0(n241), .S0(n250), .D1(n255), .S1(n240), .D2(n252), 
        .S2(n236), .D3(n238), .S3(n257), .Z(n5238) );
  HS65_LL_AOI212X4 U9710 ( .A(n265), .B(n5240), .C(n237), .D(n4927), .E(n5241), 
        .Z(n5237) );
  HS65_LL_NAND4ABX3 U9711 ( .A(n8494), .B(n8495), .C(n8496), .D(n8497), .Z(
        n3001) );
  HS65_LL_AOI212X4 U9712 ( .A(n341), .B(n8498), .C(n324), .D(n8343), .E(n8499), 
        .Z(n8497) );
  HS65_LL_MX41X7 U9713 ( .D0(n343), .S0(n330), .D1(n328), .S1(n356), .D2(n353), 
        .S2(n329), .D3(n327), .S3(n7761), .Z(n8495) );
  HS65_LL_MX41X7 U9714 ( .D0(n333), .S0(n348), .D1(n325), .S1(n347), .D2(n323), 
        .S2(n344), .D3(n355), .S3(n326), .Z(n8494) );
  HS65_LL_NAND4ABX3 U9715 ( .A(n8752), .B(n8753), .C(n8754), .D(n8755), .Z(
        n2801) );
  HS65_LL_AOI212X4 U9716 ( .A(n131), .B(n8756), .C(n111), .D(n7928), .E(n8757), 
        .Z(n8755) );
  HS65_LL_MX41X7 U9717 ( .D0(n99), .S0(n123), .D1(n119), .S1(n110), .D2(n112), 
        .S2(n122), .D3(n134), .S3(n113), .Z(n8752) );
  HS65_LL_MX41X7 U9718 ( .D0(n105), .S0(n132), .D1(n107), .S1(n136), .D2(n135), 
        .S2(n108), .D3(n106), .S3(n7738), .Z(n8753) );
  HS65_LLS_XOR2X6 U9719 ( .A(n2804), .B(n2780), .Z(n7535) );
  HS65_LLS_XOR2X6 U9720 ( .A(n2666), .B(n2897), .Z(n2706) );
  HS65_LL_NAND4ABX3 U9721 ( .A(n4285), .B(n4286), .C(n4287), .D(n4288), .Z(
        n2718) );
  HS65_LL_MX41X7 U9722 ( .D0(n437), .S0(n416), .D1(n432), .S1(n409), .D2(n411), 
        .S2(n438), .D3(n417), .S3(n3190), .Z(n4286) );
  HS65_LL_NOR4ABX2 U9723 ( .A(n3188), .B(n3845), .C(n4289), .D(n3859), .Z(
        n4288) );
  HS65_LL_MX41X7 U9724 ( .D0(n419), .S0(n436), .D1(n420), .S1(n440), .D2(n415), 
        .S2(n431), .D3(n405), .S3(n441), .Z(n4285) );
  HS65_LLS_XOR2X6 U9725 ( .A(n3209), .B(n2766), .Z(n4410) );
  HS65_LLS_XNOR2X6 U9726 ( .A(n2713), .B(n2663), .Z(n2669) );
  HS65_LLS_XOR2X6 U9727 ( .A(n2814), .B(n2790), .Z(n4378) );
  HS65_LLS_XOR2X6 U9728 ( .A(n2798), .B(n2774), .Z(n2623) );
  HS65_LLS_XOR2X6 U9729 ( .A(n2815), .B(n229), .Z(n4372) );
  HS65_LLS_XOR2X6 U9730 ( .A(n2807), .B(n51), .Z(n5965) );
  HS65_LL_NAND4ABX3 U9731 ( .A(n4226), .B(n4227), .C(n4228), .D(n4229), .Z(
        n2672) );
  HS65_LL_MX41X7 U9732 ( .D0(n637), .S0(n653), .D1(n638), .S1(n649), .D2(n633), 
        .S2(n644), .D3(n624), .S3(n650), .Z(n4226) );
  HS65_LL_MX41X7 U9733 ( .D0(n654), .S0(n634), .D1(n645), .S1(n628), .D2(n629), 
        .S2(n655), .D3(n635), .S3(n3163), .Z(n4227) );
  HS65_LL_NOR4ABX2 U9734 ( .A(n3161), .B(n3730), .C(n4230), .D(n3744), .Z(
        n4229) );
  HS65_LLS_XNOR2X6 U9735 ( .A(n2631), .B(n2637), .Z(n2685) );
  HS65_LL_NAND4ABX3 U9736 ( .A(n6943), .B(n6944), .C(n6945), .D(n6946), .Z(
        n2809) );
  HS65_LL_MX41X7 U9737 ( .D0(n276), .S0(n306), .D1(n301), .S1(n277), .D2(n300), 
        .S2(n274), .D3(n275), .S3(n6377), .Z(n6944) );
  HS65_LL_AOI212X4 U9738 ( .A(n307), .B(n6947), .C(n279), .D(n6573), .E(n6948), 
        .Z(n6946) );
  HS65_LL_MX41X7 U9739 ( .D0(n283), .S0(n292), .D1(n297), .S1(n282), .D2(n294), 
        .S2(n278), .D3(n280), .S3(n299), .Z(n6943) );
  HS65_LL_NAND4ABX3 U9740 ( .A(n3771), .B(n3772), .C(n3773), .D(n3774), .Z(
        n2703) );
  HS65_LL_MX41X7 U9741 ( .D0(n430), .S0(n413), .D1(n412), .S1(n442), .D2(n443), 
        .S2(n409), .D3(n411), .S3(n3190), .Z(n3772) );
  HS65_LL_AOI212X4 U9742 ( .A(n429), .B(n3775), .C(n407), .D(n3384), .E(n410), 
        .Z(n3774) );
  HS65_LL_MX41X7 U9743 ( .D0(n415), .S0(n431), .D1(n408), .S1(n435), .D2(n405), 
        .S2(n432), .D3(n441), .S3(n406), .Z(n3771) );
  HS65_LLS_XOR2X6 U9744 ( .A(n2808), .B(n2784), .Z(n5962) );
  HS65_LLS_XOR2X6 U9745 ( .A(n2816), .B(n2792), .Z(n4369) );
  HS65_LLS_XOR2X6 U9746 ( .A(n2799), .B(n574), .Z(n2618) );
  HS65_LLS_XNOR2X6 U9747 ( .A(n3007), .B(n2759), .Z(n6000) );
  HS65_LLS_XNOR2X6 U9748 ( .A(n3210), .B(n2767), .Z(n4407) );
  HS65_LLS_XOR2X6 U9749 ( .A(n2800), .B(n2776), .Z(n7555) );
  HS65_LLS_XNOR2X6 U9750 ( .A(n2708), .B(n2659), .Z(n2665) );
  HS65_LL_IVX9 U9751 ( .A(n2860), .Z(n197) );
  HS65_LL_IVX9 U9752 ( .A(n2882), .Z(n629) );
  HS65_LL_IVX9 U9753 ( .A(n7851), .Z(n375) );
  HS65_LL_IVX9 U9754 ( .A(n2918), .Z(n152) );
  HS65_LL_NOR4ABX2 U9755 ( .A(n7757), .B(n7758), .C(n7759), .D(n7760), .Z(
        n2898) );
  HS65_LL_MX41X7 U9756 ( .D0(n317), .S0(n351), .D1(n354), .S1(n322), .D2(n333), 
        .S2(n348), .D3(n323), .S3(n355), .Z(n7759) );
  HS65_LL_MX41X7 U9757 ( .D0(n350), .S0(n335), .D1(n329), .S1(n344), .D2(n327), 
        .S2(n352), .D3(n334), .S3(n7761), .Z(n7760) );
  HS65_LL_NOR4ABX2 U9758 ( .A(n7762), .B(n7763), .C(n7764), .D(n7765), .Z(
        n7758) );
  HS65_LL_NAND4ABX3 U9759 ( .A(n5351), .B(n5352), .C(n5353), .D(n5354), .Z(
        n2817) );
  HS65_LL_MX41X7 U9760 ( .D0(n451), .S0(n481), .D1(n476), .S1(n452), .D2(n475), 
        .S2(n449), .D3(n450), .S3(n4784), .Z(n5352) );
  HS65_LL_AOI212X4 U9761 ( .A(n482), .B(n5355), .C(n454), .D(n4980), .E(n5356), 
        .Z(n5354) );
  HS65_LL_MX41X7 U9762 ( .D0(n458), .S0(n467), .D1(n472), .S1(n457), .D2(n469), 
        .S2(n453), .D3(n455), .S3(n474), .Z(n5351) );
  HS65_LL_AOI222X2 U9763 ( .A(n639), .B(n646), .C(n661), .D(n631), .E(n640), 
        .F(n645), .Z(n4245) );
  HS65_LL_NAND4ABX3 U9764 ( .A(n3537), .B(n3538), .C(n3539), .D(n3540), .Z(
        n2652) );
  HS65_LL_MX41X7 U9765 ( .D0(n175), .S0(n153), .D1(n154), .S1(n164), .D2(n163), 
        .S2(n151), .D3(n152), .S3(n3040), .Z(n3538) );
  HS65_LL_MX41X7 U9766 ( .D0(n147), .S0(n179), .D1(n157), .S1(n177), .D2(n156), 
        .S2(n180), .D3(n158), .S3(n166), .Z(n3537) );
  HS65_LL_AOI212X4 U9767 ( .A(n173), .B(n3541), .C(n155), .D(n3257), .E(n3542), 
        .Z(n3540) );
  HS65_LL_NOR4ABX2 U9768 ( .A(n3413), .B(n3414), .C(n3415), .D(n3416), .Z(
        n2733) );
  HS65_LL_MX41X7 U9769 ( .D0(n211), .S0(n198), .D1(n199), .S1(n219), .D2(n218), 
        .S2(n196), .D3(n197), .S3(n2963), .Z(n3416) );
  HS65_LL_MX41X7 U9770 ( .D0(n192), .S0(n225), .D1(n202), .S1(n223), .D2(n201), 
        .S2(n226), .D3(n221), .S3(n203), .Z(n3415) );
  HS65_LL_AOI212X4 U9771 ( .A(n210), .B(n3417), .C(n200), .D(n3101), .E(n3418), 
        .Z(n3414) );
  HS65_LL_NAND3X5 U9772 ( .A(n7914), .B(n7915), .C(n7916), .Z(n7648) );
  HS65_LL_NOR3AX2 U9773 ( .A(n7922), .B(n7923), .C(n7924), .Z(n7915) );
  HS65_LL_NOR3AX2 U9774 ( .A(n7925), .B(n7926), .C(n7927), .Z(n7914) );
  HS65_LL_AOI212X4 U9775 ( .A(n134), .B(n100), .C(n120), .D(n98), .E(n7917), 
        .Z(n7916) );
  HS65_LL_AOI222X2 U9776 ( .A(n881), .B(n909), .C(n893), .D(n913), .E(n895), 
        .F(n908), .Z(n2564) );
  HS65_LL_NAND3X5 U9777 ( .A(n1403), .B(n1404), .C(n1405), .Z(n1125) );
  HS65_LL_NOR3AX2 U9778 ( .A(n1230), .B(n1357), .C(n1335), .Z(n1404) );
  HS65_LL_NOR3X4 U9779 ( .A(n1275), .B(n1409), .C(n1315), .Z(n1403) );
  HS65_LL_AOI212X4 U9780 ( .A(n844), .B(n873), .C(n863), .D(n839), .E(n1406), 
        .Z(n1405) );
  HS65_LL_NAND3X5 U9781 ( .A(n2155), .B(n2156), .C(n2157), .Z(n1877) );
  HS65_LL_NOR3AX2 U9782 ( .A(n1982), .B(n2109), .C(n2087), .Z(n2156) );
  HS65_LL_NOR3X4 U9783 ( .A(n2027), .B(n2161), .C(n2067), .Z(n2155) );
  HS65_LL_AOI212X4 U9784 ( .A(n762), .B(n791), .C(n781), .D(n757), .E(n2158), 
        .Z(n2157) );
  HS65_LL_NAND3X5 U9785 ( .A(n1779), .B(n1780), .C(n1781), .Z(n1501) );
  HS65_LL_NOR3AX2 U9786 ( .A(n1606), .B(n1733), .C(n1711), .Z(n1780) );
  HS65_LL_NOR3X4 U9787 ( .A(n1651), .B(n1785), .C(n1691), .Z(n1779) );
  HS65_LL_AOI212X4 U9788 ( .A(n803), .B(n832), .C(n822), .D(n798), .E(n1782), 
        .Z(n1781) );
  HS65_LL_NAND3X5 U9789 ( .A(n4174), .B(n4175), .C(n4176), .Z(n3919) );
  HS65_LL_NOR3X4 U9790 ( .A(n3530), .B(n3093), .C(n3508), .Z(n4175) );
  HS65_LL_NOR3X4 U9791 ( .A(n4180), .B(n3487), .C(n3433), .Z(n4174) );
  HS65_LL_AOI212X4 U9792 ( .A(n221), .B(n194), .C(n193), .D(n224), .E(n4177), 
        .Z(n4176) );
  HS65_LL_NAND3X5 U9793 ( .A(n4026), .B(n4027), .C(n4028), .Z(n2850) );
  HS65_LL_NOR3AX2 U9794 ( .A(n3377), .B(n3884), .C(n3862), .Z(n4027) );
  HS65_LL_NOR3X4 U9795 ( .A(n4032), .B(n3843), .C(n3791), .Z(n4026) );
  HS65_LL_AOI212X4 U9796 ( .A(n441), .B(n417), .C(n418), .D(n433), .E(n4029), 
        .Z(n4028) );
  HS65_LL_NOR4ABX2 U9797 ( .A(n8662), .B(n8663), .C(n8664), .D(n8665), .Z(
        n2777) );
  HS65_LL_MX41X7 U9798 ( .D0(n579), .S0(n603), .D1(n599), .S1(n590), .D2(n592), 
        .S2(n602), .D3(n614), .S3(n593), .Z(n8664) );
  HS65_LL_MX41X7 U9799 ( .D0(n585), .S0(n612), .D1(n587), .S1(n616), .D2(n615), 
        .S2(n588), .D3(n586), .S3(n7700), .Z(n8665) );
  HS65_LL_AOI212X4 U9800 ( .A(n611), .B(n8666), .C(n591), .D(n7830), .E(n8667), 
        .Z(n8663) );
  HS65_LL_AOI212X4 U9801 ( .A(n335), .B(n346), .C(n328), .D(n340), .E(n8628), 
        .Z(n8627) );
  HS65_LL_CB4I6X9 U9802 ( .A(n324), .B(n327), .C(n347), .D(n8521), .Z(n8628)
         );
  HS65_LL_NAND3X5 U9803 ( .A(n8901), .B(n8902), .C(n8903), .Z(n8623) );
  HS65_LL_NOR3X4 U9804 ( .A(n8593), .B(n8337), .C(n8570), .Z(n8902) );
  HS65_LL_NOR3X4 U9805 ( .A(n8909), .B(n8553), .C(n8609), .Z(n8901) );
  HS65_LL_AOI212X4 U9806 ( .A(n355), .B(n334), .C(n332), .D(n345), .E(n8904), 
        .Z(n8903) );
  HS65_LL_IVX9 U9807 ( .A(n2246), .Z(n896) );
  HS65_LL_IVX9 U9808 ( .A(n1118), .Z(n855) );
  HS65_LL_IVX9 U9809 ( .A(n1494), .Z(n814) );
  HS65_LL_IVX9 U9810 ( .A(n1870), .Z(n773) );
  HS65_LL_AOI212X4 U9811 ( .A(n368), .B(n385), .C(n376), .D(n389), .E(n8656), 
        .Z(n8655) );
  HS65_LL_CB4I6X9 U9812 ( .A(n371), .B(n375), .C(n386), .D(n8306), .Z(n8656)
         );
  HS65_LL_AOI222X2 U9813 ( .A(n888), .B(n909), .C(n885), .D(n2287), .E(n916), 
        .F(n895), .Z(n2487) );
  HS65_LL_AOI222X2 U9814 ( .A(n765), .B(n786), .C(n762), .D(n1911), .E(n793), 
        .F(n772), .Z(n2111) );
  HS65_LL_AOI222X2 U9815 ( .A(n847), .B(n868), .C(n844), .D(n1159), .E(n875), 
        .F(n854), .Z(n1359) );
  HS65_LL_AOI222X2 U9816 ( .A(n806), .B(n827), .C(n803), .D(n1535), .E(n834), 
        .F(n813), .Z(n1735) );
  HS65_LL_AOI222X2 U9817 ( .A(n400), .B(n365), .C(n393), .D(n372), .E(n373), 
        .F(n389), .Z(n8645) );
  HS65_LL_AOI212X4 U9818 ( .A(n634), .B(n647), .C(n630), .D(n659), .E(n4279), 
        .Z(n4274) );
  HS65_LL_CB4I6X9 U9819 ( .A(n626), .B(n629), .C(n648), .D(n3687), .Z(n4279)
         );
  HS65_LLS_XNOR2X6 U9820 ( .A(n2810), .B(n5940), .Z(n6016) );
  HS65_LLS_XNOR2X6 U9821 ( .A(n2818), .B(n4347), .Z(n4423) );
  HS65_LLS_XOR2X6 U9822 ( .A(n2774), .B(n7532), .Z(n7640) );
  HS65_LLS_XOR2X6 U9823 ( .A(n2802), .B(n7532), .Z(n7605) );
  HS65_LL_NOR4ABX2 U9824 ( .A(n4044), .B(n4045), .C(n4046), .D(n4047), .Z(
        n2745) );
  HS65_LL_MX41X7 U9825 ( .D0(n215), .S0(n195), .D1(n226), .S1(n196), .D2(n197), 
        .S2(n214), .D3(n194), .S3(n2963), .Z(n4047) );
  HS65_LL_MX41X7 U9826 ( .D0(n191), .S0(n216), .D1(n188), .S1(n220), .D2(n192), 
        .S2(n225), .D3(n201), .S3(n221), .Z(n4046) );
  HS65_LL_NOR4ABX2 U9827 ( .A(n2961), .B(n3490), .C(n4048), .D(n3505), .Z(
        n4045) );
  HS65_LLS_XOR2X6 U9828 ( .A(n3000), .B(n7546), .Z(n7549) );
  HS65_LL_NOR4ABX2 U9829 ( .A(n4141), .B(n4142), .C(n4143), .D(n4144), .Z(
        n4095) );
  HS65_LL_NAND4ABX3 U9830 ( .A(n3593), .B(n3651), .C(n2920), .D(n3610), .Z(
        n4143) );
  HS65_LL_NAND4ABX3 U9831 ( .A(n3581), .B(n3259), .C(n3051), .D(n3558), .Z(
        n4144) );
  HS65_LL_NOR3AX2 U9832 ( .A(n4149), .B(n3570), .C(n3283), .Z(n4142) );
  HS65_LL_NOR4ABX2 U9833 ( .A(n4107), .B(n4108), .C(n4109), .D(n4110), .Z(
        n4080) );
  HS65_LL_NAND3X5 U9834 ( .A(n3559), .B(n3247), .C(n3576), .Z(n4110) );
  HS65_LL_NAND4ABX3 U9835 ( .A(n3649), .B(n3037), .C(n3614), .D(n3639), .Z(
        n4109) );
  HS65_LL_AOI222X2 U9836 ( .A(n142), .B(n178), .C(n158), .D(n164), .E(n156), 
        .F(n172), .Z(n4107) );
  HS65_LL_NOR4ABX2 U9837 ( .A(n4273), .B(n4274), .C(n4275), .D(n4276), .Z(
        n2877) );
  HS65_LL_NAND4ABX3 U9838 ( .A(n3156), .B(n3325), .C(n3673), .D(n3749), .Z(
        n4275) );
  HS65_LL_NAND3AX6 U9839 ( .A(n3727), .B(n3768), .C(n3663), .Z(n4276) );
  HS65_LL_AOI222X2 U9840 ( .A(n638), .B(n646), .C(n651), .D(n625), .E(n658), 
        .F(n624), .Z(n4273) );
  HS65_LL_NOR4ABX2 U9841 ( .A(n1469), .B(n1470), .C(n1471), .D(n1472), .Z(
        n1131) );
  HS65_LL_NAND4ABX3 U9842 ( .A(n1192), .B(n1232), .C(n1273), .D(n1337), .Z(
        n1471) );
  HS65_LL_NOR3AX2 U9843 ( .A(n1356), .B(n1262), .C(n1314), .Z(n1470) );
  HS65_LL_AOI222X2 U9844 ( .A(n868), .B(n839), .C(n854), .D(n874), .E(n847), 
        .F(n860), .Z(n1469) );
  HS65_LL_NOR4ABX2 U9845 ( .A(n2221), .B(n2222), .C(n2223), .D(n2224), .Z(
        n1883) );
  HS65_LL_NAND4ABX3 U9846 ( .A(n1944), .B(n1984), .C(n2025), .D(n2089), .Z(
        n2223) );
  HS65_LL_NOR3AX2 U9847 ( .A(n2108), .B(n2014), .C(n2066), .Z(n2222) );
  HS65_LL_AOI222X2 U9848 ( .A(n786), .B(n757), .C(n772), .D(n792), .E(n765), 
        .F(n778), .Z(n2221) );
  HS65_LL_NOR4ABX2 U9849 ( .A(n2597), .B(n2598), .C(n2599), .D(n2600), .Z(
        n2259) );
  HS65_LL_NAND4ABX3 U9850 ( .A(n2320), .B(n2360), .C(n2401), .D(n2465), .Z(
        n2599) );
  HS65_LL_NOR3AX2 U9851 ( .A(n2484), .B(n2390), .C(n2442), .Z(n2598) );
  HS65_LL_AOI222X2 U9852 ( .A(n909), .B(n880), .C(n895), .D(n915), .E(n888), 
        .F(n901), .Z(n2597) );
  HS65_LL_NOR4ABX2 U9853 ( .A(n1845), .B(n1846), .C(n1847), .D(n1848), .Z(
        n1507) );
  HS65_LL_NAND4ABX3 U9854 ( .A(n1568), .B(n1608), .C(n1649), .D(n1713), .Z(
        n1847) );
  HS65_LL_NOR3AX2 U9855 ( .A(n1732), .B(n1638), .C(n1690), .Z(n1846) );
  HS65_LL_AOI222X2 U9856 ( .A(n827), .B(n798), .C(n813), .D(n833), .E(n806), 
        .F(n819), .Z(n1845) );
  HS65_LL_NOR4ABX2 U9857 ( .A(n4332), .B(n4333), .C(n4334), .D(n4335), .Z(
        n2847) );
  HS65_LL_NAND4ABX3 U9858 ( .A(n3182), .B(n3379), .C(n3788), .D(n3864), .Z(
        n4334) );
  HS65_LL_NOR3AX2 U9859 ( .A(n3883), .B(n3779), .C(n3842), .Z(n4333) );
  HS65_LL_AOI222X2 U9860 ( .A(n420), .B(n433), .C(n442), .D(n406), .E(n427), 
        .F(n405), .Z(n4332) );
  HS65_LL_NOR4ABX2 U9861 ( .A(n8951), .B(n8952), .C(n8953), .D(n8954), .Z(
        n8491) );
  HS65_LL_NAND4ABX3 U9862 ( .A(n7989), .B(n8218), .C(n8257), .D(n8108), .Z(
        n8954) );
  HS65_LL_NAND4ABX3 U9863 ( .A(n8090), .B(n8305), .C(n8955), .D(n8078), .Z(
        n8953) );
  HS65_LL_AOI222X2 U9864 ( .A(n395), .B(n366), .C(n375), .D(n399), .E(n374), 
        .F(n396), .Z(n8951) );
  HS65_LL_NOR4ABX2 U9865 ( .A(n8891), .B(n8892), .C(n8893), .D(n8894), .Z(
        n8869) );
  HS65_LL_NAND4ABX3 U9866 ( .A(n8059), .B(n8605), .C(n8559), .D(n8341), .Z(
        n8894) );
  HS65_LL_NAND4ABX3 U9867 ( .A(n8322), .B(n8519), .C(n8895), .D(n8354), .Z(
        n8893) );
  HS65_LL_AOI222X2 U9868 ( .A(n353), .B(n322), .C(n327), .D(n350), .E(n325), 
        .F(n356), .Z(n8891) );
  HS65_LL_NAND4ABX3 U9869 ( .A(n4254), .B(n4255), .C(n4256), .D(n4257), .Z(
        n3948) );
  HS65_LL_AOI222X2 U9870 ( .A(n653), .B(n639), .C(n650), .D(n625), .E(n624), 
        .F(n659), .Z(n4256) );
  HS65_LL_NAND4ABX3 U9871 ( .A(n3345), .B(n3710), .C(n3690), .D(n3319), .Z(
        n4255) );
  HS65_LL_NAND4ABX3 U9872 ( .A(n3153), .B(n3700), .C(n3722), .D(n3740), .Z(
        n4254) );
  HS65_LL_NAND4ABX3 U9873 ( .A(n4313), .B(n4314), .C(n4315), .D(n4316), .Z(
        n3968) );
  HS65_LL_NAND4ABX3 U9874 ( .A(n3399), .B(n3825), .C(n3805), .D(n3373), .Z(
        n4314) );
  HS65_LL_NAND4ABX3 U9875 ( .A(n3179), .B(n3840), .C(n3817), .D(n3855), .Z(
        n4313) );
  HS65_LL_AOI222X2 U9876 ( .A(n436), .B(n421), .C(n441), .D(n406), .E(n405), 
        .F(n428), .Z(n4315) );
  HS65_LL_NAND3X5 U9877 ( .A(n4003), .B(n4004), .C(n4005), .Z(n2880) );
  HS65_LL_NOR3AX2 U9878 ( .A(n3323), .B(n3769), .C(n3747), .Z(n4004) );
  HS65_LL_NOR3X4 U9879 ( .A(n4009), .B(n3728), .C(n3676), .Z(n4003) );
  HS65_LL_AOI212X4 U9880 ( .A(n650), .B(n635), .C(n636), .D(n646), .E(n4006), 
        .Z(n4005) );
  HS65_LL_NAND4ABX3 U9881 ( .A(n1428), .B(n1429), .C(n1430), .D(n1431), .Z(
        n1402) );
  HS65_LL_MX41X7 U9882 ( .D0(n842), .S0(n871), .D1(n847), .S1(n866), .D2(n863), 
        .S2(n840), .D3(n852), .S3(n864), .Z(n1428) );
  HS65_LL_NAND3AX6 U9883 ( .A(n1238), .B(n1342), .C(n1449), .Z(n1429) );
  HS65_LL_AOI212X4 U9884 ( .A(n844), .B(n1285), .C(n870), .D(n849), .E(n1432), 
        .Z(n1431) );
  HS65_LL_NAND4ABX3 U9885 ( .A(n2180), .B(n2181), .C(n2182), .D(n2183), .Z(
        n2154) );
  HS65_LL_MX41X7 U9886 ( .D0(n760), .S0(n789), .D1(n765), .S1(n784), .D2(n781), 
        .S2(n758), .D3(n770), .S3(n782), .Z(n2180) );
  HS65_LL_NAND3AX6 U9887 ( .A(n1990), .B(n2094), .C(n2201), .Z(n2181) );
  HS65_LL_AOI212X4 U9888 ( .A(n762), .B(n2037), .C(n788), .D(n767), .E(n2184), 
        .Z(n2183) );
  HS65_LL_NAND4ABX3 U9889 ( .A(n1804), .B(n1805), .C(n1806), .D(n1807), .Z(
        n1778) );
  HS65_LL_MX41X7 U9890 ( .D0(n801), .S0(n830), .D1(n806), .S1(n825), .D2(n822), 
        .S2(n799), .D3(n811), .S3(n823), .Z(n1804) );
  HS65_LL_NAND3AX6 U9891 ( .A(n1614), .B(n1718), .C(n1825), .Z(n1805) );
  HS65_LL_AOI212X4 U9892 ( .A(n803), .B(n1661), .C(n829), .D(n808), .E(n1808), 
        .Z(n1807) );
  HS65_LL_NAND4ABX3 U9893 ( .A(n2556), .B(n2557), .C(n2558), .D(n2559), .Z(
        n2530) );
  HS65_LL_AOI212X4 U9894 ( .A(n885), .B(n2413), .C(n911), .D(n890), .E(n2560), 
        .Z(n2559) );
  HS65_LL_MX41X7 U9895 ( .D0(n883), .S0(n912), .D1(n888), .S1(n907), .D2(n904), 
        .S2(n881), .D3(n893), .S3(n905), .Z(n2556) );
  HS65_LL_NAND3AX6 U9896 ( .A(n2366), .B(n2470), .C(n2577), .Z(n2557) );
  HS65_LL_NAND4ABX3 U9897 ( .A(n4052), .B(n4053), .C(n4054), .D(n4055), .Z(
        n3920) );
  HS65_LL_MX41X7 U9898 ( .D0(n211), .S0(n200), .D1(n209), .S1(n198), .D2(n193), 
        .S2(n218), .D3(n215), .S3(n191), .Z(n4052) );
  HS65_LL_NAND3AX6 U9899 ( .A(n3102), .B(n3515), .C(n4065), .Z(n4053) );
  HS65_LL_AOI212X4 U9900 ( .A(n221), .B(n3461), .C(n199), .D(n220), .E(n4056), 
        .Z(n4055) );
  HS65_LL_NAND4ABX3 U9901 ( .A(n4232), .B(n4233), .C(n4234), .D(n4235), .Z(
        n4002) );
  HS65_LL_AOI212X4 U9902 ( .A(n650), .B(n3703), .C(n630), .D(n649), .E(n4236), 
        .Z(n4235) );
  HS65_LL_MX41X7 U9903 ( .D0(n661), .S0(n626), .D1(n658), .S1(n631), .D2(n636), 
        .S2(n652), .D3(n654), .S3(n637), .Z(n4232) );
  HS65_LL_NAND3AX6 U9904 ( .A(n3331), .B(n3754), .C(n4253), .Z(n4233) );
  HS65_LL_NAND4ABX3 U9905 ( .A(n4291), .B(n4292), .C(n4293), .D(n4294), .Z(
        n4025) );
  HS65_LL_MX41X7 U9906 ( .D0(n430), .S0(n407), .D1(n427), .S1(n413), .D2(n418), 
        .S2(n443), .D3(n437), .S3(n419), .Z(n4291) );
  HS65_LL_NAND3AX6 U9907 ( .A(n3385), .B(n3869), .C(n4312), .Z(n4292) );
  HS65_LL_AOI212X4 U9908 ( .A(n441), .B(n3818), .C(n412), .D(n440), .E(n4295), 
        .Z(n4294) );
  HS65_LL_NAND3X5 U9909 ( .A(n7185), .B(n7186), .C(n7187), .Z(n6045) );
  HS65_LL_AND3X9 U9910 ( .A(n6511), .B(n6881), .C(n6895), .Z(n7186) );
  HS65_LL_NOR3X4 U9911 ( .A(n7191), .B(n6861), .C(n6942), .Z(n7185) );
  HS65_LL_AOI212X4 U9912 ( .A(n56), .B(n76), .C(n88), .D(n55), .E(n7188), .Z(
        n7187) );
  HS65_LL_NAND3X5 U9913 ( .A(n8961), .B(n8962), .C(n8963), .Z(n8637) );
  HS65_LL_NOR3X4 U9914 ( .A(n8291), .B(n8104), .C(n8269), .Z(n8962) );
  HS65_LL_NOR3X4 U9915 ( .A(n8969), .B(n8250), .C(n8224), .Z(n8961) );
  HS65_LL_AOI212X4 U9916 ( .A(n393), .B(n370), .C(n369), .D(n384), .E(n8964), 
        .Z(n8963) );
  HS65_LLS_XNOR2X6 U9917 ( .A(n2815), .B(n7), .Z(n4434) );
  HS65_LL_NAND4ABX3 U9918 ( .A(n6598), .B(n6599), .C(n6600), .D(n6601), .Z(
        n6069) );
  HS65_LL_NAND4ABX3 U9919 ( .A(n6662), .B(n6663), .C(n6664), .D(n6665), .Z(
        n6599) );
  HS65_LL_MX41X7 U9920 ( .D0(n537), .S0(n553), .D1(n561), .S1(n546), .D2(n533), 
        .S2(n552), .D3(n542), .S3(n550), .Z(n6598) );
  HS65_LL_AOI212X4 U9921 ( .A(n555), .B(n6602), .C(n538), .D(n560), .E(n6603), 
        .Z(n6601) );
  HS65_LL_NAND4ABX3 U9922 ( .A(n6719), .B(n6720), .C(n6721), .D(n6722), .Z(
        n6125) );
  HS65_LL_NAND4ABX3 U9923 ( .A(n6783), .B(n6784), .C(n6785), .D(n6786), .Z(
        n6720) );
  HS65_LL_MX41X7 U9924 ( .D0(n494), .S0(n510), .D1(n503), .S1(n518), .D2(n492), 
        .S2(n509), .D3(n499), .S3(n507), .Z(n6719) );
  HS65_LL_AOI212X4 U9925 ( .A(n512), .B(n6723), .C(n495), .D(n517), .E(n6724), 
        .Z(n6722) );
  HS65_LL_NAND4ABX3 U9926 ( .A(n5005), .B(n5006), .C(n5007), .D(n5008), .Z(
        n4476) );
  HS65_LL_NAND4ABX3 U9927 ( .A(n5069), .B(n5070), .C(n5071), .D(n5072), .Z(
        n5006) );
  HS65_LL_MX41X7 U9928 ( .D0(n15), .S0(n31), .D1(n39), .S1(n24), .D2(n11), 
        .S2(n30), .D3(n20), .S3(n28), .Z(n5005) );
  HS65_LL_AOI212X4 U9929 ( .A(n33), .B(n5009), .C(n16), .D(n38), .E(n5010), 
        .Z(n5008) );
  HS65_LL_NAND4ABX3 U9930 ( .A(n5127), .B(n5128), .C(n5129), .D(n5130), .Z(
        n4532) );
  HS65_LL_NAND4ABX3 U9931 ( .A(n5191), .B(n5192), .C(n5193), .D(n5194), .Z(
        n5128) );
  HS65_LL_MX41X7 U9932 ( .D0(n670), .S0(n686), .D1(n679), .S1(n694), .D2(n668), 
        .S2(n685), .D3(n675), .S3(n683), .Z(n5127) );
  HS65_LL_AOI212X4 U9933 ( .A(n688), .B(n5131), .C(n671), .D(n693), .E(n5132), 
        .Z(n5130) );
  HS65_LL_NAND4ABX3 U9934 ( .A(n6837), .B(n6838), .C(n6839), .D(n6840), .Z(
        n6178) );
  HS65_LL_NAND4ABX3 U9935 ( .A(n6899), .B(n6900), .C(n6901), .D(n6902), .Z(
        n6838) );
  HS65_LL_MX41X7 U9936 ( .D0(n55), .S0(n74), .D1(n63), .S1(n82), .D2(n67), 
        .S2(n77), .D3(n60), .S3(n72), .Z(n6837) );
  HS65_LL_AOI212X4 U9937 ( .A(n76), .B(n6841), .C(n54), .D(n80), .E(n6842), 
        .Z(n6840) );
  HS65_LL_NAND4ABX3 U9938 ( .A(n5245), .B(n5246), .C(n5247), .D(n5248), .Z(
        n4585) );
  HS65_LL_NAND4ABX3 U9939 ( .A(n5307), .B(n5308), .C(n5309), .D(n5310), .Z(
        n5246) );
  HS65_LL_MX41X7 U9940 ( .D0(n244), .S0(n256), .D1(n234), .S1(n268), .D2(n246), 
        .S2(n259), .D3(n238), .S3(n254), .Z(n5245) );
  HS65_LL_AOI212X4 U9941 ( .A(n257), .B(n5249), .C(n242), .D(n266), .E(n5250), 
        .Z(n5248) );
  HS65_LL_NAND4ABX3 U9942 ( .A(n5360), .B(n5361), .C(n5362), .D(n5363), .Z(
        n4602) );
  HS65_LL_NAND4ABX3 U9943 ( .A(n5422), .B(n5423), .C(n5424), .D(n5425), .Z(
        n5361) );
  HS65_LL_MX41X7 U9944 ( .D0(n461), .S0(n473), .D1(n451), .S1(n485), .D2(n463), 
        .S2(n476), .D3(n455), .S3(n471), .Z(n5360) );
  HS65_LL_AOI212X4 U9945 ( .A(n474), .B(n5364), .C(n459), .D(n483), .E(n5365), 
        .Z(n5363) );
  HS65_LL_NAND4ABX3 U9946 ( .A(n6952), .B(n6953), .C(n6954), .D(n6955), .Z(
        n6195) );
  HS65_LL_NAND4ABX3 U9947 ( .A(n7014), .B(n7015), .C(n7016), .D(n7017), .Z(
        n6953) );
  HS65_LL_MX41X7 U9948 ( .D0(n286), .S0(n298), .D1(n276), .S1(n310), .D2(n288), 
        .S2(n301), .D3(n280), .S3(n296), .Z(n6952) );
  HS65_LL_AOI212X4 U9949 ( .A(n299), .B(n6956), .C(n284), .D(n308), .E(n6957), 
        .Z(n6955) );
  HS65_LL_NAND4ABX3 U9950 ( .A(n8670), .B(n8671), .C(n8672), .D(n8673), .Z(
        n8002) );
  HS65_LL_NAND4ABX3 U9951 ( .A(n8716), .B(n8717), .C(n8718), .D(n7797), .Z(
        n8671) );
  HS65_LL_MX41X7 U9952 ( .D0(n578), .S0(n617), .D1(n585), .S1(n609), .D2(n582), 
        .S2(n616), .D3(n593), .S3(n598), .Z(n8670) );
  HS65_LL_AOI212X4 U9953 ( .A(n614), .B(n8674), .C(n576), .D(n608), .E(n8675), 
        .Z(n8673) );
  HS65_LL_NAND4ABX3 U9954 ( .A(n8760), .B(n8761), .C(n8762), .D(n8763), .Z(
        n8015) );
  HS65_LL_NAND4ABX3 U9955 ( .A(n8806), .B(n8807), .C(n8808), .D(n7896), .Z(
        n8761) );
  HS65_LL_MX41X7 U9956 ( .D0(n98), .S0(n137), .D1(n105), .S1(n129), .D2(n102), 
        .S2(n136), .D3(n113), .S3(n118), .Z(n8760) );
  HS65_LL_AOI212X4 U9957 ( .A(n134), .B(n8764), .C(n96), .D(n128), .E(n8765), 
        .Z(n8763) );
  HS65_LL_NOR4ABX2 U9958 ( .A(n8956), .B(n8957), .C(n8958), .D(n8959), .Z(
        n8636) );
  HS65_LL_NAND4ABX3 U9959 ( .A(n8113), .B(n7991), .C(n8249), .D(n8210), .Z(
        n8959) );
  HS65_LL_NAND4ABX3 U9960 ( .A(n8077), .B(n8307), .C(n8960), .D(n8227), .Z(
        n8958) );
  HS65_LL_AOI222X2 U9961 ( .A(n384), .B(n365), .C(n392), .D(n378), .E(n363), 
        .F(n383), .Z(n8956) );
  HS65_LL_NAND4ABX3 U9962 ( .A(n5272), .B(n5273), .C(n5274), .D(n5275), .Z(
        n4909) );
  HS65_LL_NAND3X5 U9963 ( .A(n5284), .B(n5285), .C(n5286), .Z(n5273) );
  HS65_LL_NOR4ABX2 U9964 ( .A(n5276), .B(n5277), .C(n5278), .D(n5279), .Z(
        n5275) );
  HS65_LL_NAND4ABX3 U9965 ( .A(n5287), .B(n5288), .C(n5289), .D(n5290), .Z(
        n5272) );
  HS65_LL_NAND4ABX3 U9966 ( .A(n6864), .B(n6865), .C(n6866), .D(n6867), .Z(
        n6502) );
  HS65_LL_NAND3X5 U9967 ( .A(n6876), .B(n6877), .C(n6878), .Z(n6865) );
  HS65_LL_NOR4ABX2 U9968 ( .A(n6868), .B(n6869), .C(n6870), .D(n6871), .Z(
        n6867) );
  HS65_LL_NAND4ABX3 U9969 ( .A(n6879), .B(n6880), .C(n6881), .D(n6882), .Z(
        n6864) );
  HS65_LL_NAND4ABX3 U9970 ( .A(n6979), .B(n6980), .C(n6981), .D(n6982), .Z(
        n6555) );
  HS65_LL_NAND3X5 U9971 ( .A(n6991), .B(n6992), .C(n6993), .Z(n6980) );
  HS65_LL_NOR4ABX2 U9972 ( .A(n6983), .B(n6984), .C(n6985), .D(n6986), .Z(
        n6982) );
  HS65_LL_NAND4ABX3 U9973 ( .A(n6994), .B(n6995), .C(n6996), .D(n6997), .Z(
        n6979) );
  HS65_LL_NOR4ABX2 U9974 ( .A(n5925), .B(n5926), .C(n5927), .D(n5928), .Z(
        n4510) );
  HS65_LL_NAND4ABX3 U9975 ( .A(n4945), .B(n5461), .C(n5447), .D(n5932), .Z(
        n5927) );
  HS65_LL_AOI222X2 U9976 ( .A(n470), .B(n463), .C(n451), .D(n481), .E(n464), 
        .F(n469), .Z(n5925) );
  HS65_LL_NAND4X9 U9977 ( .A(n4984), .B(n4779), .C(n5372), .D(n5436), .Z(n5928) );
  HS65_LL_NOR4ABX2 U9978 ( .A(n7517), .B(n7518), .C(n7519), .D(n7520), .Z(
        n6103) );
  HS65_LL_NAND4ABX3 U9979 ( .A(n6538), .B(n7053), .C(n7039), .D(n7524), .Z(
        n7519) );
  HS65_LL_AOI222X2 U9980 ( .A(n295), .B(n288), .C(n276), .D(n306), .E(n289), 
        .F(n294), .Z(n7517) );
  HS65_LL_NAND4X9 U9981 ( .A(n6577), .B(n6372), .C(n6964), .D(n7028), .Z(n7520) );
  HS65_LL_NOR4ABX2 U9982 ( .A(n5866), .B(n5867), .C(n5868), .D(n5869), .Z(
        n4449) );
  HS65_LL_NAND4ABX3 U9983 ( .A(n4892), .B(n5346), .C(n5332), .D(n5873), .Z(
        n5868) );
  HS65_LL_AOI222X2 U9984 ( .A(n253), .B(n246), .C(n234), .D(n264), .E(n247), 
        .F(n252), .Z(n5866) );
  HS65_LL_NAND4X9 U9985 ( .A(n4931), .B(n4752), .C(n5257), .D(n5321), .Z(n5869) );
  HS65_LL_NOR4ABX2 U9986 ( .A(n7462), .B(n7463), .C(n7464), .D(n7465), .Z(
        n6042) );
  HS65_LL_NAND4ABX3 U9987 ( .A(n6485), .B(n6938), .C(n6924), .D(n7467), .Z(
        n7464) );
  HS65_LL_AOI222X2 U9988 ( .A(n88), .B(n67), .C(n63), .D(n78), .E(n68), .F(n89), .Z(n7462) );
  HS65_LL_NAND4X9 U9989 ( .A(n6524), .B(n6333), .C(n6849), .D(n6913), .Z(n7465) );
  HS65_LL_NOR4ABX2 U9990 ( .A(n5762), .B(n5763), .C(n5764), .D(n5765), .Z(
        n5687) );
  HS65_LL_NAND4ABX3 U9991 ( .A(n4817), .B(n5231), .C(n5216), .D(n5766), .Z(
        n5764) );
  HS65_LL_AOI222X2 U9992 ( .A(n700), .B(n668), .C(n679), .D(n697), .E(n666), 
        .F(n702), .Z(n5762) );
  HS65_LL_NAND4X9 U9993 ( .A(n4858), .B(n4633), .C(n5140), .D(n5205), .Z(n5765) );
  HS65_LL_NOR4ABX2 U9994 ( .A(n7354), .B(n7355), .C(n7356), .D(n7357), .Z(
        n7279) );
  HS65_LL_NAND4ABX3 U9995 ( .A(n6410), .B(n6823), .C(n6808), .D(n7358), .Z(
        n7356) );
  HS65_LL_AOI222X2 U9996 ( .A(n524), .B(n492), .C(n503), .D(n521), .E(n490), 
        .F(n526), .Z(n7354) );
  HS65_LL_NAND4X9 U9997 ( .A(n6451), .B(n6226), .C(n6732), .D(n6797), .Z(n7357) );
  HS65_LL_NOR4ABX2 U9998 ( .A(n6646), .B(n6647), .C(n6648), .D(n6649), .Z(
        n6264) );
  HS65_LL_NAND3AX6 U9999 ( .A(n6650), .B(n6651), .C(n6652), .Z(n6648) );
  HS65_LL_MX41X7 U10000 ( .D0(n531), .S0(n553), .D1(n563), .S1(n533), .D2(n564), .S2(n538), .D3(n551), .S3(n536), .Z(n6649) );
  HS65_LL_NOR4ABX2 U10001 ( .A(n6658), .B(n6659), .C(n6660), .D(n6661), .Z(
        n6646) );
  HS65_LL_NOR4ABX2 U10002 ( .A(n5053), .B(n5054), .C(n5055), .D(n5056), .Z(
        n4671) );
  HS65_LL_NAND3AX6 U10003 ( .A(n5057), .B(n5058), .C(n5059), .Z(n5055) );
  HS65_LL_MX41X7 U10004 ( .D0(n9), .S0(n31), .D1(n41), .S1(n11), .D2(n42), 
        .S2(n16), .D3(n29), .S3(n14), .Z(n5056) );
  HS65_LL_NOR4ABX2 U10005 ( .A(n5065), .B(n5066), .C(n5067), .D(n5068), .Z(
        n5053) );
  HS65_LL_NOR4ABX2 U10006 ( .A(n6767), .B(n6768), .C(n6769), .D(n6770), .Z(
        n6403) );
  HS65_LL_NAND3AX6 U10007 ( .A(n6771), .B(n6772), .C(n6773), .Z(n6769) );
  HS65_LL_MX41X7 U10008 ( .D0(n489), .S0(n510), .D1(n492), .S1(n520), .D2(n521), .S2(n495), .D3(n508), .S3(n493), .Z(n6770) );
  HS65_LL_NOR4ABX2 U10009 ( .A(n6779), .B(n6780), .C(n6781), .D(n6782), .Z(
        n6767) );
  HS65_LL_NOR4ABX2 U10010 ( .A(n5175), .B(n5176), .C(n5177), .D(n5178), .Z(
        n4810) );
  HS65_LL_NAND3AX6 U10011 ( .A(n5179), .B(n5180), .C(n5181), .Z(n5177) );
  HS65_LL_MX41X7 U10012 ( .D0(n665), .S0(n686), .D1(n668), .S1(n696), .D2(n697), .S2(n671), .D3(n684), .S3(n669), .Z(n5178) );
  HS65_LL_NOR4ABX2 U10013 ( .A(n5187), .B(n5188), .C(n5189), .D(n5190), .Z(
        n5175) );
  HS65_LL_NOR4ABX2 U10014 ( .A(n6883), .B(n6884), .C(n6885), .D(n6886), .Z(
        n6478) );
  HS65_LL_NAND3AX6 U10015 ( .A(n6887), .B(n6888), .C(n6889), .Z(n6885) );
  HS65_LL_MX41X7 U10016 ( .D0(n69), .S0(n74), .D1(n67), .S1(n81), .D2(n78), 
        .S2(n54), .D3(n73), .S3(n57), .Z(n6886) );
  HS65_LL_NOR4ABX2 U10017 ( .A(n6895), .B(n6896), .C(n6897), .D(n6898), .Z(
        n6883) );
  HS65_LL_NOR4ABX2 U10018 ( .A(n5291), .B(n5292), .C(n5293), .D(n5294), .Z(
        n4885) );
  HS65_LL_NAND3AX6 U10019 ( .A(n5295), .B(n5296), .C(n5297), .Z(n5293) );
  HS65_LL_MX41X7 U10020 ( .D0(n245), .S0(n256), .D1(n246), .S1(n267), .D2(n264), .S2(n242), .D3(n258), .S3(n241), .Z(n5294) );
  HS65_LL_NOR4ABX2 U10021 ( .A(n5303), .B(n5304), .C(n5305), .D(n5306), .Z(
        n5291) );
  HS65_LL_NOR4ABX2 U10022 ( .A(n5406), .B(n5407), .C(n5408), .D(n5409), .Z(
        n4938) );
  HS65_LL_NAND3AX6 U10023 ( .A(n5410), .B(n5411), .C(n5412), .Z(n5408) );
  HS65_LL_MX41X7 U10024 ( .D0(n462), .S0(n473), .D1(n463), .S1(n484), .D2(n481), .S2(n459), .D3(n475), .S3(n458), .Z(n5409) );
  HS65_LL_NOR4ABX2 U10025 ( .A(n5418), .B(n5419), .C(n5420), .D(n5421), .Z(
        n5406) );
  HS65_LL_NOR4ABX2 U10026 ( .A(n6998), .B(n6999), .C(n7000), .D(n7001), .Z(
        n6531) );
  HS65_LL_NAND3AX6 U10027 ( .A(n7002), .B(n7003), .C(n7004), .Z(n7000) );
  HS65_LL_MX41X7 U10028 ( .D0(n287), .S0(n298), .D1(n288), .S1(n309), .D2(n306), .S2(n284), .D3(n300), .S3(n283), .Z(n7001) );
  HS65_LL_NOR4ABX2 U10029 ( .A(n7010), .B(n7011), .C(n7012), .D(n7013), .Z(
        n6998) );
  HS65_LL_NOR4ABX2 U10030 ( .A(n4169), .B(n4170), .C(n4171), .D(n4172), .Z(
        n4057) );
  HS65_LL_NAND4ABX3 U10031 ( .A(n3486), .B(n2955), .C(n3105), .D(n3459), .Z(
        n4172) );
  HS65_LL_NAND4ABX3 U10032 ( .A(n3122), .B(n3444), .C(n4173), .D(n3430), .Z(
        n4171) );
  HS65_LL_AOI222X2 U10033 ( .A(n190), .B(n224), .C(n211), .D(n198), .E(n189), 
        .F(n226), .Z(n4169) );
  HS65_LL_NOR4ABX2 U10034 ( .A(n3640), .B(n3641), .C(n3642), .D(n3643), .Z(
        n3226) );
  HS65_LL_MX41X7 U10035 ( .D0(n142), .S0(n165), .D1(n145), .S1(n174), .D2(n175), .S2(n150), .D3(n147), .S3(n163), .Z(n3643) );
  HS65_LL_NAND4ABX3 U10036 ( .A(n3644), .B(n3645), .C(n3646), .D(n3647), .Z(
        n3642) );
  HS65_LL_NOR3AX2 U10037 ( .A(n3648), .B(n3649), .C(n3650), .Z(n3641) );
  HS65_LL_NOR4ABX2 U10038 ( .A(n8896), .B(n8897), .C(n8898), .D(n8899), .Z(
        n8621) );
  HS65_LL_NAND4ABX3 U10039 ( .A(n8346), .B(n8060), .C(n8551), .D(n8513), .Z(
        n8899) );
  HS65_LL_NAND4ABX3 U10040 ( .A(n8353), .B(n8520), .C(n8900), .D(n8608), .Z(
        n8898) );
  HS65_LL_AOI222X2 U10041 ( .A(n345), .B(n319), .C(n343), .D(n330), .E(n320), 
        .F(n344), .Z(n8896) );
  HS65_LL_NOR4ABX2 U10042 ( .A(n7784), .B(n7785), .C(n7786), .D(n7787), .Z(
        n7695) );
  HS65_LL_NAND4ABX3 U10043 ( .A(n7788), .B(n7789), .C(n7790), .D(n7791), .Z(
        n7787) );
  HS65_LL_NAND4ABX3 U10044 ( .A(n7792), .B(n7793), .C(n7794), .D(n7795), .Z(
        n7786) );
  HS65_LL_AOI222X2 U10045 ( .A(n600), .B(n582), .C(n585), .D(n612), .E(n583), 
        .F(n602), .Z(n7784) );
  HS65_LL_NOR4ABX2 U10046 ( .A(n7883), .B(n7884), .C(n7885), .D(n7886), .Z(
        n7733) );
  HS65_LL_NAND4ABX3 U10047 ( .A(n7887), .B(n7888), .C(n7889), .D(n7890), .Z(
        n7886) );
  HS65_LL_NAND4ABX3 U10048 ( .A(n7891), .B(n7892), .C(n7893), .D(n7894), .Z(
        n7885) );
  HS65_LL_AOI222X2 U10049 ( .A(n120), .B(n102), .C(n105), .D(n132), .E(n103), 
        .F(n122), .Z(n7883) );
  HS65_LL_NOR4ABX2 U10050 ( .A(n7292), .B(n7293), .C(n7294), .D(n7295), .Z(
        n7249) );
  HS65_LL_NAND4ABX3 U10051 ( .A(n6613), .B(n6148), .C(n6314), .D(n6676), .Z(
        n7295) );
  HS65_LL_NAND4ABX3 U10052 ( .A(n6272), .B(n6701), .C(n7296), .D(n6686), .Z(
        n7294) );
  HS65_LL_AOI222X2 U10053 ( .A(n533), .B(n567), .C(n546), .D(n564), .E(n532), 
        .F(n569), .Z(n7292) );
  HS65_LL_NOR4ABX2 U10054 ( .A(n5700), .B(n5701), .C(n5702), .D(n5703), .Z(
        n5657) );
  HS65_LL_NAND4ABX3 U10055 ( .A(n5020), .B(n4555), .C(n4721), .D(n5083), .Z(
        n5703) );
  HS65_LL_NAND4ABX3 U10056 ( .A(n4679), .B(n5108), .C(n5704), .D(n5093), .Z(
        n5702) );
  HS65_LL_AOI222X2 U10057 ( .A(n11), .B(n45), .C(n24), .D(n42), .E(n10), .F(
        n47), .Z(n5700) );
  HS65_LL_NOR4ABX2 U10058 ( .A(n2471), .B(n2472), .C(n2473), .D(n2474), .Z(
        n2337) );
  HS65_LL_NAND3X5 U10059 ( .A(n2475), .B(n2476), .C(n2477), .Z(n2473) );
  HS65_LL_MX41X7 U10060 ( .D0(n909), .S0(n890), .D1(n892), .S1(n903), .D2(n883), .S2(n910), .D3(n881), .S3(n906), .Z(n2474) );
  HS65_LL_NOR4ABX2 U10061 ( .A(n2479), .B(n2480), .C(n2481), .D(n2482), .Z(
        n2472) );
  HS65_LL_NOR4ABX2 U10062 ( .A(n1343), .B(n1344), .C(n1345), .D(n1346), .Z(
        n1209) );
  HS65_LL_NAND3X5 U10063 ( .A(n1347), .B(n1348), .C(n1349), .Z(n1345) );
  HS65_LL_MX41X7 U10064 ( .D0(n868), .S0(n849), .D1(n851), .S1(n862), .D2(n842), .S2(n869), .D3(n840), .S3(n865), .Z(n1346) );
  HS65_LL_NOR4ABX2 U10065 ( .A(n1351), .B(n1352), .C(n1353), .D(n1354), .Z(
        n1344) );
  HS65_LL_NOR4ABX2 U10066 ( .A(n2095), .B(n2096), .C(n2097), .D(n2098), .Z(
        n1961) );
  HS65_LL_NAND3X5 U10067 ( .A(n2099), .B(n2100), .C(n2101), .Z(n2097) );
  HS65_LL_MX41X7 U10068 ( .D0(n786), .S0(n767), .D1(n769), .S1(n780), .D2(n760), .S2(n787), .D3(n758), .S3(n783), .Z(n2098) );
  HS65_LL_NOR4ABX2 U10069 ( .A(n2103), .B(n2104), .C(n2105), .D(n2106), .Z(
        n2096) );
  HS65_LL_NOR4ABX2 U10070 ( .A(n1719), .B(n1720), .C(n1721), .D(n1722), .Z(
        n1585) );
  HS65_LL_NAND3X5 U10071 ( .A(n1723), .B(n1724), .C(n1725), .Z(n1721) );
  HS65_LL_MX41X7 U10072 ( .D0(n827), .S0(n808), .D1(n810), .S1(n821), .D2(n801), .S2(n828), .D3(n799), .S3(n824), .Z(n1722) );
  HS65_LL_NOR4ABX2 U10073 ( .A(n1727), .B(n1728), .C(n1729), .D(n1730), .Z(
        n1720) );
  HS65_LL_NOR4ABX2 U10074 ( .A(n3755), .B(n3756), .C(n3757), .D(n3758), .Z(
        n3301) );
  HS65_LL_MX41X7 U10075 ( .D0(n638), .S0(n649), .D1(n659), .S1(n639), .D2(n661), .S2(n634), .D3(n652), .S3(n633), .Z(n3758) );
  HS65_LL_NAND3X5 U10076 ( .A(n3759), .B(n3760), .C(n3761), .Z(n3757) );
  HS65_LL_NOR4ABX2 U10077 ( .A(n3767), .B(n3768), .C(n3769), .D(n3770), .Z(
        n3755) );
  HS65_LL_NOR4ABX2 U10078 ( .A(n3870), .B(n3871), .C(n3872), .D(n3873), .Z(
        n3355) );
  HS65_LL_MX41X7 U10079 ( .D0(n420), .S0(n440), .D1(n428), .S1(n421), .D2(n430), .S2(n416), .D3(n443), .S3(n415), .Z(n3873) );
  HS65_LL_NAND3X5 U10080 ( .A(n3874), .B(n3875), .C(n3876), .Z(n3872) );
  HS65_LL_NOR4ABX2 U10081 ( .A(n3878), .B(n3879), .C(n3880), .D(n3881), .Z(
        n3871) );
  HS65_LL_NOR4ABX2 U10082 ( .A(n3516), .B(n3517), .C(n3518), .D(n3519), .Z(
        n3070) );
  HS65_LL_NAND3X5 U10083 ( .A(n3520), .B(n3521), .C(n3522), .Z(n3518) );
  HS65_LL_MX41X7 U10084 ( .D0(n188), .S0(n220), .D1(n212), .S1(n190), .D2(n211), .S2(n195), .D3(n218), .S3(n192), .Z(n3519) );
  HS65_LL_NOR4ABX2 U10085 ( .A(n3524), .B(n3525), .C(n3526), .D(n3527), .Z(
        n3517) );
  HS65_LL_NOR4ABX2 U10086 ( .A(n8704), .B(n8705), .C(n8706), .D(n8707), .Z(
        n8375) );
  HS65_LL_MX41X7 U10087 ( .D0(n584), .S0(n617), .D1(n582), .S1(n610), .D2(n612), .S2(n576), .D3(n615), .S3(n579), .Z(n8707) );
  HS65_LL_NAND3X5 U10088 ( .A(n8708), .B(n7810), .C(n8709), .Z(n8706) );
  HS65_LL_NOR4ABX2 U10089 ( .A(n8713), .B(n7824), .C(n8714), .D(n8715), .Z(
        n8704) );
  HS65_LL_NOR4ABX2 U10090 ( .A(n8794), .B(n8795), .C(n8796), .D(n8797), .Z(
        n8427) );
  HS65_LL_MX41X7 U10091 ( .D0(n104), .S0(n137), .D1(n102), .S1(n130), .D2(n132), .S2(n96), .D3(n135), .S3(n99), .Z(n8797) );
  HS65_LL_NAND3X5 U10092 ( .A(n8798), .B(n7908), .C(n8799), .Z(n8796) );
  HS65_LL_NOR4ABX2 U10093 ( .A(n8803), .B(n7922), .C(n8804), .D(n8805), .Z(
        n8794) );
  HS65_LL_NOR4ABX2 U10094 ( .A(n8277), .B(n8278), .C(n8279), .D(n8280), .Z(
        n8068) );
  HS65_LL_MX41X7 U10095 ( .D0(n394), .S0(n366), .D1(n389), .S1(n365), .D2(n392), .S2(n368), .D3(n367), .S3(n395), .Z(n8280) );
  HS65_LL_NAND3X5 U10096 ( .A(n8281), .B(n8282), .C(n8283), .Z(n8279) );
  HS65_LL_NOR4ABX2 U10097 ( .A(n8285), .B(n8286), .C(n8287), .D(n8288), .Z(
        n8278) );
  HS65_LL_NAND4ABX3 U10098 ( .A(n3303), .B(n3304), .C(n3305), .D(n3306), .Z(
        n3145) );
  HS65_LL_NAND4ABX3 U10099 ( .A(n3332), .B(n3333), .C(n3334), .D(n3335), .Z(
        n3304) );
  HS65_LL_NOR4ABX2 U10100 ( .A(n3307), .B(n3308), .C(n3309), .D(n3310), .Z(
        n3306) );
  HS65_LL_MX41X7 U10101 ( .D0(n637), .S0(n655), .D1(n640), .S1(n661), .D2(n624), .S2(n648), .D3(n629), .S3(n658), .Z(n3303) );
  HS65_LL_NOR4ABX2 U10102 ( .A(n8579), .B(n8580), .C(n8581), .D(n8582), .Z(
        n8314) );
  HS65_LL_MX41X7 U10103 ( .D0(n354), .S0(n322), .D1(n340), .S1(n319), .D2(n343), .S2(n335), .D3(n333), .S3(n353), .Z(n8582) );
  HS65_LL_NAND3AX6 U10104 ( .A(n8583), .B(n8584), .C(n8585), .Z(n8581) );
  HS65_LL_NOR4ABX2 U10105 ( .A(n8587), .B(n8588), .C(n8589), .D(n8590), .Z(
        n8580) );
  HS65_LL_NAND4ABX3 U10106 ( .A(n3357), .B(n3358), .C(n3359), .D(n3360), .Z(
        n3171) );
  HS65_LL_NAND4ABX3 U10107 ( .A(n3386), .B(n3387), .C(n3388), .D(n3389), .Z(
        n3358) );
  HS65_LL_NOR4ABX2 U10108 ( .A(n3361), .B(n3362), .C(n3363), .D(n3364), .Z(
        n3360) );
  HS65_LL_MX41X7 U10109 ( .D0(n419), .S0(n438), .D1(n422), .S1(n430), .D2(n405), .S2(n435), .D3(n411), .S3(n427), .Z(n3357) );
  HS65_LL_OAI31X5 U10110 ( .A(n883), .B(n886), .C(n885), .D(n903), .Z(n2342)
         );
  HS65_LL_OAI31X5 U10111 ( .A(n760), .B(n763), .C(n762), .D(n780), .Z(n1966)
         );
  HS65_LL_NAND4ABX3 U10112 ( .A(n8743), .B(n8744), .C(n8745), .D(n8746), .Z(
        n8139) );
  HS65_LL_AOI222X2 U10113 ( .A(n609), .B(n579), .C(n591), .D(n617), .E(n578), 
        .F(n611), .Z(n8745) );
  HS65_LL_AOI212X4 U10114 ( .A(n600), .B(n7684), .C(n604), .D(n8747), .E(n8748), .Z(n8746) );
  HS65_LL_NAND4ABX3 U10115 ( .A(n8749), .B(n8750), .C(n7791), .D(n8751), .Z(
        n8744) );
  HS65_LL_OAI31X5 U10116 ( .A(n842), .B(n845), .C(n844), .D(n862), .Z(n1214)
         );
  HS65_LL_OAI31X5 U10117 ( .A(n801), .B(n804), .C(n803), .D(n821), .Z(n1590)
         );
  HS65_LL_NOR3X4 U10118 ( .A(n7800), .B(n7628), .C(n7680), .Z(n7780) );
  HS65_LL_IVX9 U10119 ( .A(n1486), .Z(n831) );
  HS65_LL_IVX9 U10120 ( .A(n2238), .Z(n913) );
  HS65_LL_IVX9 U10121 ( .A(n1110), .Z(n872) );
  HS65_LL_IVX9 U10122 ( .A(n1862), .Z(n790) );
  HS65_LL_NOR3X4 U10123 ( .A(n4450), .B(n4451), .C(n4452), .Z(n4444) );
  HS65_LL_NOR3X4 U10124 ( .A(n5490), .B(n5675), .C(n5569), .Z(n5759) );
  HS65_LL_NOR3X4 U10125 ( .A(n7082), .B(n7267), .C(n7161), .Z(n7351) );
  HS65_LL_NOR3X4 U10126 ( .A(n6043), .B(n6044), .C(n6045), .Z(n6037) );
  HS65_LL_NOR3X4 U10127 ( .A(n7755), .B(n8485), .C(n8637), .Z(n8633) );
  HS65_LL_NOR3X4 U10128 ( .A(n3910), .B(n4088), .C(n3986), .Z(n4104) );
  HS65_LL_NOR3X4 U10129 ( .A(n5476), .B(n5645), .C(n5505), .Z(n5697) );
  HS65_LL_NOR3X4 U10130 ( .A(n7068), .B(n7237), .C(n7097), .Z(n7289) );
  HS65_LL_NAND4ABX3 U10131 ( .A(n4243), .B(n4244), .C(n4245), .D(n4246), .Z(
        n2879) );
  HS65_LL_NAND4ABX3 U10132 ( .A(n3333), .B(n3155), .C(n3726), .D(n3702), .Z(
        n4244) );
  HS65_LL_NAND4ABX3 U10133 ( .A(n3349), .B(n3675), .C(n3685), .D(n4247), .Z(
        n4243) );
  HS65_LL_NOR4ABX2 U10134 ( .A(n3767), .B(n3712), .C(n3324), .D(n3748), .Z(
        n4246) );
  HS65_LL_NAND4ABX3 U10135 ( .A(n4302), .B(n4303), .C(n4304), .D(n4305), .Z(
        n2849) );
  HS65_LL_AOI222X2 U10136 ( .A(n421), .B(n433), .C(n430), .D(n413), .E(n422), 
        .F(n432), .Z(n4304) );
  HS65_LL_NAND4ABX3 U10137 ( .A(n3841), .B(n3181), .C(n3388), .D(n3816), .Z(
        n4303) );
  HS65_LL_NAND4ABX3 U10138 ( .A(n3403), .B(n3790), .C(n3800), .D(n4306), .Z(
        n4302) );
  HS65_LL_NAND2X7 U10139 ( .A(n392), .B(n362), .Z(n8210) );
  HS65_LLS_XNOR2X6 U10140 ( .A(n3008), .B(n272), .Z(n5956) );
  HS65_LLS_XNOR2X6 U10141 ( .A(n3211), .B(n447), .Z(n4363) );
  HS65_LL_NAND4ABX3 U10142 ( .A(n4238), .B(n4239), .C(n4240), .D(n4241), .Z(
        n3940) );
  HS65_LL_AOI222X2 U10143 ( .A(n652), .B(n638), .C(n654), .D(n629), .E(n651), 
        .F(n627), .Z(n4240) );
  HS65_LL_NAND4ABX3 U10144 ( .A(n3686), .B(n3705), .C(n3674), .D(n4242), .Z(
        n4238) );
  HS65_LL_NAND4ABX3 U10145 ( .A(n3348), .B(n3309), .C(n3154), .D(n3322), .Z(
        n4239) );
  HS65_LL_NOR4ABX2 U10146 ( .A(n8879), .B(n8880), .C(n8881), .D(n8882), .Z(
        n7772) );
  HS65_LL_NAND3AX6 U10147 ( .A(n8610), .B(n8591), .C(n8883), .Z(n8882) );
  HS65_LL_MX41X7 U10148 ( .D0(n324), .S0(n343), .D1(n342), .S1(n330), .D2(n353), .S2(n332), .D3(n317), .S3(n350), .Z(n8881) );
  HS65_LL_AOI212X4 U10149 ( .A(n355), .B(n8507), .C(n328), .D(n354), .E(n8884), 
        .Z(n8880) );
  HS65_LL_NOR3X4 U10150 ( .A(n3312), .B(n3313), .C(n2979), .Z(n3305) );
  HS65_LL_NOR3X4 U10151 ( .A(n2347), .B(n2348), .C(n2269), .Z(n2340) );
  HS65_LL_NOR3X4 U10152 ( .A(n1971), .B(n1972), .C(n1893), .Z(n1964) );
  HS65_LL_NOR3X4 U10153 ( .A(n1219), .B(n1220), .C(n1141), .Z(n1212) );
  HS65_LL_NOR3X4 U10154 ( .A(n1595), .B(n1596), .C(n1517), .Z(n1588) );
  HS65_LL_NOR3X4 U10155 ( .A(n3366), .B(n3367), .C(n2990), .Z(n3359) );
  HS65_LL_NOR4ABX2 U10156 ( .A(n8939), .B(n8940), .C(n8941), .D(n8942), .Z(
        n7754) );
  HS65_LL_NAND3X5 U10157 ( .A(n8289), .B(n8226), .C(n8943), .Z(n8942) );
  HS65_LL_MX41X7 U10158 ( .D0(n371), .S0(n392), .D1(n390), .S1(n378), .D2(n395), .S2(n369), .D3(n362), .S3(n399), .Z(n8941) );
  HS65_LL_AOI212X4 U10159 ( .A(n393), .B(n8204), .C(n376), .D(n394), .E(n8944), 
        .Z(n8940) );
  HS65_LL_NOR4ABX2 U10160 ( .A(n8530), .B(n8531), .C(n8532), .D(n8533), .Z(
        n7944) );
  HS65_LL_NAND4ABX3 U10161 ( .A(n8534), .B(n8535), .C(n8536), .D(n8537), .Z(
        n8533) );
  HS65_LL_MX41X7 U10162 ( .D0(n332), .S0(n354), .D1(n342), .S1(n330), .D2(n356), .S2(n319), .D3(n326), .S3(n346), .Z(n8532) );
  HS65_LL_AOI212X4 U10163 ( .A(n355), .B(n8538), .C(n335), .D(n339), .E(n8539), 
        .Z(n8531) );
  HS65_LL_NOR2X6 U10164 ( .A(n390), .B(n389), .Z(n8240) );
  HS65_LL_NAND4ABX3 U10165 ( .A(n7251), .B(n7252), .C(n7253), .D(n7254), .Z(
        n7069) );
  HS65_LL_NAND4ABX3 U10166 ( .A(n534), .B(n6688), .C(n6612), .D(n6294), .Z(
        n7252) );
  HS65_LL_AOI222X2 U10167 ( .A(n531), .B(n551), .C(n545), .D(n559), .E(n543), 
        .F(n552), .Z(n7253) );
  HS65_LL_NAND4ABX3 U10168 ( .A(n6271), .B(n6312), .C(n6702), .D(n7255), .Z(
        n7251) );
  HS65_LL_NAND4ABX3 U10169 ( .A(n5659), .B(n5660), .C(n5661), .D(n5662), .Z(
        n5477) );
  HS65_LL_NAND4ABX3 U10170 ( .A(n12), .B(n5095), .C(n5019), .D(n4701), .Z(
        n5660) );
  HS65_LL_AOI222X2 U10171 ( .A(n9), .B(n29), .C(n23), .D(n37), .E(n21), .F(n30), .Z(n5661) );
  HS65_LL_NAND4ABX3 U10172 ( .A(n4678), .B(n4719), .C(n5109), .D(n5663), .Z(
        n5659) );
  HS65_LL_NOR2X6 U10173 ( .A(n435), .B(n443), .Z(n3973) );
  HS65_LL_NOR2X6 U10174 ( .A(n648), .B(n652), .Z(n3935) );
  HS65_LL_NOR2X6 U10175 ( .A(n658), .B(n659), .Z(n3717) );
  HS65_LL_NAND2X7 U10176 ( .A(n395), .B(n362), .Z(n8257) );
  HS65_LL_NAND4ABX3 U10177 ( .A(n5906), .B(n5907), .C(n5908), .D(n5909), .Z(
        n5557) );
  HS65_LL_AOI222X2 U10178 ( .A(n462), .B(n475), .C(n450), .D(n478), .E(n457), 
        .F(n476), .Z(n5908) );
  HS65_LL_NAND4ABX3 U10179 ( .A(n4778), .B(n5375), .C(n5459), .D(n4967), .Z(
        n5907) );
  HS65_LL_NOR4ABX2 U10180 ( .A(n5425), .B(n5414), .C(n5434), .D(n5394), .Z(
        n5909) );
  HS65_LL_NAND4ABX3 U10181 ( .A(n7498), .B(n7499), .C(n7500), .D(n7501), .Z(
        n7149) );
  HS65_LL_AOI222X2 U10182 ( .A(n287), .B(n300), .C(n275), .D(n303), .E(n282), 
        .F(n301), .Z(n7500) );
  HS65_LL_NAND4ABX3 U10183 ( .A(n6371), .B(n6967), .C(n7051), .D(n6560), .Z(
        n7499) );
  HS65_LL_NOR4ABX2 U10184 ( .A(n7017), .B(n7006), .C(n7026), .D(n6986), .Z(
        n7501) );
  HS65_LL_NAND4ABX3 U10185 ( .A(n5847), .B(n5848), .C(n5849), .D(n5850), .Z(
        n5535) );
  HS65_LL_AOI222X2 U10186 ( .A(n245), .B(n258), .C(n233), .D(n261), .E(n240), 
        .F(n259), .Z(n5849) );
  HS65_LL_NAND4ABX3 U10187 ( .A(n4751), .B(n5260), .C(n5344), .D(n4914), .Z(
        n5848) );
  HS65_LL_NOR4ABX2 U10188 ( .A(n5310), .B(n5299), .C(n5319), .D(n5279), .Z(
        n5850) );
  HS65_LL_NAND4ABX3 U10189 ( .A(n7439), .B(n7440), .C(n7441), .D(n7442), .Z(
        n7127) );
  HS65_LL_AOI222X2 U10190 ( .A(n69), .B(n73), .C(n64), .D(n85), .E(n62), .F(
        n77), .Z(n7441) );
  HS65_LL_NAND4ABX3 U10191 ( .A(n6332), .B(n6852), .C(n6936), .D(n6507), .Z(
        n7440) );
  HS65_LL_NOR4ABX2 U10192 ( .A(n6902), .B(n6891), .C(n6911), .D(n6871), .Z(
        n7442) );
  HS65_LL_NOR2X6 U10193 ( .A(n888), .B(n892), .Z(n2432) );
  HS65_LL_NOR2X6 U10194 ( .A(n765), .B(n769), .Z(n2056) );
  HS65_LL_NOR2X6 U10195 ( .A(n847), .B(n851), .Z(n1304) );
  HS65_LL_NOR2X6 U10196 ( .A(n806), .B(n810), .Z(n1680) );
  HS65_LL_NOR4ABX2 U10197 ( .A(n8858), .B(n8859), .C(n8860), .D(n8861), .Z(
        n7771) );
  HS65_LL_NAND4ABX3 U10198 ( .A(n8361), .B(n8333), .C(n8536), .D(n8524), .Z(
        n8861) );
  HS65_LL_NAND4ABX3 U10199 ( .A(n8511), .B(n8550), .C(n8565), .D(n8054), .Z(
        n8860) );
  HS65_LL_AOI222X2 U10200 ( .A(n351), .B(n319), .C(n355), .D(n326), .E(n323), 
        .F(n340), .Z(n8858) );
  HS65_LL_NOR2X6 U10201 ( .A(n347), .B(n353), .Z(n8629) );
  HS65_LL_NOR4ABX2 U10202 ( .A(n8645), .B(n8646), .C(n8647), .D(n8648), .Z(
        n7753) );
  HS65_LL_NAND4ABX3 U10203 ( .A(n8076), .B(n8100), .C(n8234), .D(n8299), .Z(
        n8648) );
  HS65_LL_NAND4ABX3 U10204 ( .A(n8208), .B(n8248), .C(n8263), .D(n7986), .Z(
        n8647) );
  HS65_LL_NOR4ABX2 U10205 ( .A(n8650), .B(n8115), .C(n8288), .D(n8222), .Z(
        n8646) );
  HS65_LL_NAND4ABX3 U10206 ( .A(n2033), .B(n2034), .C(n2035), .D(n2036), .Z(
        n1922) );
  HS65_LL_AOI212X4 U10207 ( .A(n757), .B(n2037), .C(n759), .D(n2038), .E(n2039), .Z(n2036) );
  HS65_LL_MX41X7 U10208 ( .D0(n784), .S0(n771), .D1(n772), .S1(n792), .D2(n770), .S2(n782), .D3(n760), .S3(n779), .Z(n2033) );
  HS65_LL_AOI222X2 U10209 ( .A(n783), .B(n765), .C(n789), .D(n767), .E(n781), 
        .F(n773), .Z(n2035) );
  HS65_LL_NAND4ABX3 U10210 ( .A(n1281), .B(n1282), .C(n1283), .D(n1284), .Z(
        n1170) );
  HS65_LL_AOI212X4 U10211 ( .A(n839), .B(n1285), .C(n841), .D(n1286), .E(n1287), .Z(n1284) );
  HS65_LL_MX41X7 U10212 ( .D0(n866), .S0(n853), .D1(n854), .S1(n874), .D2(n852), .S2(n864), .D3(n842), .S3(n861), .Z(n1281) );
  HS65_LL_AOI222X2 U10213 ( .A(n865), .B(n847), .C(n871), .D(n849), .E(n863), 
        .F(n855), .Z(n1283) );
  HS65_LL_NOR4ABX2 U10214 ( .A(n9073), .B(n9074), .C(n9075), .D(n9076), .Z(
        n7654) );
  HS65_LL_NAND4ABX3 U10215 ( .A(n8185), .B(n8805), .C(n8774), .D(n8841), .Z(
        n9076) );
  HS65_LL_MX41X7 U10216 ( .D0(n103), .S0(n137), .D1(n105), .S1(n136), .D2(n107), .S2(n129), .D3(n135), .S3(n108), .Z(n9075) );
  HS65_LL_NOR4ABX2 U10217 ( .A(n8827), .B(n109), .C(n8448), .D(n8177), .Z(
        n9073) );
  HS65_LL_NOR4ABX2 U10218 ( .A(n9015), .B(n9016), .C(n9017), .D(n9018), .Z(
        n7634) );
  HS65_LL_NAND4ABX3 U10219 ( .A(n8134), .B(n8715), .C(n8684), .D(n8751), .Z(
        n9018) );
  HS65_LL_MX41X7 U10220 ( .D0(n583), .S0(n617), .D1(n585), .S1(n616), .D2(n587), .S2(n609), .D3(n615), .S3(n588), .Z(n9017) );
  HS65_LL_NOR4ABX2 U10221 ( .A(n8737), .B(n589), .C(n8396), .D(n8154), .Z(
        n9015) );
  HS65_LL_NAND4ABX3 U10222 ( .A(n1657), .B(n1658), .C(n1659), .D(n1660), .Z(
        n1546) );
  HS65_LL_AOI212X4 U10223 ( .A(n798), .B(n1661), .C(n800), .D(n1662), .E(n1663), .Z(n1660) );
  HS65_LL_MX41X7 U10224 ( .D0(n825), .S0(n812), .D1(n813), .S1(n833), .D2(n811), .S2(n823), .D3(n801), .S3(n820), .Z(n1657) );
  HS65_LL_AOI222X2 U10225 ( .A(n824), .B(n806), .C(n830), .D(n808), .E(n822), 
        .F(n814), .Z(n1659) );
  HS65_LL_NAND4ABX3 U10226 ( .A(n2409), .B(n2410), .C(n2411), .D(n2412), .Z(
        n2298) );
  HS65_LL_AOI212X4 U10227 ( .A(n880), .B(n2413), .C(n882), .D(n2414), .E(n2415), .Z(n2412) );
  HS65_LL_MX41X7 U10228 ( .D0(n907), .S0(n894), .D1(n895), .S1(n915), .D2(n893), .S2(n905), .D3(n883), .S3(n902), .Z(n2409) );
  HS65_LL_AOI222X2 U10229 ( .A(n906), .B(n888), .C(n912), .D(n890), .E(n904), 
        .F(n896), .Z(n2411) );
  HS65_LL_NOR4ABX2 U10230 ( .A(n5894), .B(n5895), .C(n5896), .D(n5897), .Z(
        n5550) );
  HS65_LL_NAND4ABX3 U10231 ( .A(n5422), .B(n4974), .C(n4948), .D(n5442), .Z(
        n5897) );
  HS65_LL_NAND4ABX3 U10232 ( .A(n4785), .B(n5433), .C(n5396), .D(n5385), .Z(
        n5896) );
  HS65_LL_AOI222X2 U10233 ( .A(n463), .B(n477), .C(n455), .D(n474), .E(n484), 
        .F(n453), .Z(n5894) );
  HS65_LL_NOR4ABX2 U10234 ( .A(n5835), .B(n5836), .C(n5837), .D(n5838), .Z(
        n5528) );
  HS65_LL_NAND4ABX3 U10235 ( .A(n5307), .B(n4921), .C(n4895), .D(n5327), .Z(
        n5838) );
  HS65_LL_NAND4ABX3 U10236 ( .A(n4758), .B(n5318), .C(n5281), .D(n5270), .Z(
        n5837) );
  HS65_LL_AOI222X2 U10237 ( .A(n246), .B(n260), .C(n238), .D(n257), .E(n267), 
        .F(n236), .Z(n5835) );
  HS65_LL_NOR4ABX2 U10238 ( .A(n7486), .B(n7487), .C(n7488), .D(n7489), .Z(
        n7142) );
  HS65_LL_NAND4ABX3 U10239 ( .A(n7014), .B(n6567), .C(n6541), .D(n7034), .Z(
        n7489) );
  HS65_LL_NAND4ABX3 U10240 ( .A(n6378), .B(n7025), .C(n6988), .D(n6977), .Z(
        n7488) );
  HS65_LL_AOI222X2 U10241 ( .A(n288), .B(n302), .C(n280), .D(n299), .E(n309), 
        .F(n278), .Z(n7486) );
  HS65_LL_NOR4ABX2 U10242 ( .A(n5795), .B(n5796), .C(n5797), .D(n5798), .Z(
        n5674) );
  HS65_LL_NAND4ABX3 U10243 ( .A(n5191), .B(n4846), .C(n4820), .D(n5211), .Z(
        n5798) );
  HS65_LL_NAND4ABX3 U10244 ( .A(n4639), .B(n5202), .C(n5164), .D(n5153), .Z(
        n5797) );
  HS65_LL_AOI222X2 U10245 ( .A(n668), .B(n690), .C(n675), .D(n688), .E(n696), 
        .F(n674), .Z(n5795) );
  HS65_LL_NOR4ABX2 U10246 ( .A(n7387), .B(n7388), .C(n7389), .D(n7390), .Z(
        n7266) );
  HS65_LL_NAND4ABX3 U10247 ( .A(n6783), .B(n6439), .C(n6413), .D(n6803), .Z(
        n7390) );
  HS65_LL_NAND4ABX3 U10248 ( .A(n6232), .B(n6794), .C(n6756), .D(n6745), .Z(
        n7389) );
  HS65_LL_AOI222X2 U10249 ( .A(n492), .B(n514), .C(n499), .D(n512), .E(n520), 
        .F(n498), .Z(n7387) );
  HS65_LL_NOR4ABX2 U10250 ( .A(n7427), .B(n7428), .C(n7429), .D(n7430), .Z(
        n7120) );
  HS65_LL_NAND4ABX3 U10251 ( .A(n6899), .B(n6514), .C(n6488), .D(n6919), .Z(
        n7430) );
  HS65_LL_NAND4ABX3 U10252 ( .A(n6339), .B(n6910), .C(n6873), .D(n6862), .Z(
        n7429) );
  HS65_LL_AOI222X2 U10253 ( .A(n67), .B(n83), .C(n60), .D(n76), .E(n81), .F(
        n59), .Z(n7427) );
  HS65_LL_NOR4ABX2 U10254 ( .A(n5733), .B(n5734), .C(n5735), .D(n5736), .Z(
        n5644) );
  HS65_LL_NAND4ABX3 U10255 ( .A(n5069), .B(n4708), .C(n4681), .D(n5105), .Z(
        n5736) );
  HS65_LL_NAND4ABX3 U10256 ( .A(n5029), .B(n5044), .C(n5081), .D(n4562), .Z(
        n5735) );
  HS65_LL_AOI222X2 U10257 ( .A(n11), .B(n35), .C(n20), .D(n33), .E(n41), .F(
        n19), .Z(n5733) );
  HS65_LL_NOR4ABX2 U10258 ( .A(n7325), .B(n7326), .C(n7327), .D(n7328), .Z(
        n7236) );
  HS65_LL_NAND4ABX3 U10259 ( .A(n6662), .B(n6301), .C(n6274), .D(n6698), .Z(
        n7328) );
  HS65_LL_NAND4ABX3 U10260 ( .A(n6622), .B(n6637), .C(n6674), .D(n6155), .Z(
        n7327) );
  HS65_LL_AOI222X2 U10261 ( .A(n533), .B(n557), .C(n542), .D(n555), .E(n563), 
        .F(n541), .Z(n7325) );
  HS65_LL_NOR4ABX2 U10262 ( .A(n3589), .B(n3590), .C(n3591), .D(n3592), .Z(
        n2907) );
  HS65_LL_NAND4ABX3 U10263 ( .A(n3593), .B(n3594), .C(n3595), .D(n3596), .Z(
        n3592) );
  HS65_LL_MX41X7 U10264 ( .D0(n148), .S0(n165), .D1(n153), .S1(n172), .D2(n145), .S2(n164), .D3(n158), .S3(n3597), .Z(n3591) );
  HS65_LL_AOI212X4 U10265 ( .A(n166), .B(n3598), .C(n150), .D(n171), .E(n3599), 
        .Z(n3590) );
  HS65_LL_NAND4ABX3 U10266 ( .A(n4129), .B(n4130), .C(n4131), .D(n4132), .Z(
        n3988) );
  HS65_LL_NAND4ABX3 U10267 ( .A(n3258), .B(n3049), .C(n3272), .D(n3038), .Z(
        n4130) );
  HS65_LL_NOR4ABX2 U10268 ( .A(n3571), .B(n3262), .C(n3552), .D(n3587), .Z(
        n4131) );
  HS65_LL_NOR4ABX2 U10269 ( .A(n3619), .B(n3600), .C(n3655), .D(n3627), .Z(
        n4132) );
  HS65_LL_NOR4ABX2 U10270 ( .A(n3821), .B(n3822), .C(n3823), .D(n3824), .Z(
        n2987) );
  HS65_LL_NAND4ABX3 U10271 ( .A(n3825), .B(n3826), .C(n3827), .D(n3828), .Z(
        n3824) );
  HS65_LL_MX41X7 U10272 ( .D0(n418), .S0(n440), .D1(n427), .S1(n413), .D2(n442), .S2(n421), .D3(n406), .S3(n434), .Z(n3823) );
  HS65_LL_AOI212X4 U10273 ( .A(n441), .B(n3829), .C(n416), .D(n426), .E(n3830), 
        .Z(n3822) );
  HS65_LL_NOR4ABX2 U10274 ( .A(n3465), .B(n3466), .C(n3467), .D(n3468), .Z(
        n2864) );
  HS65_LL_NAND4ABX3 U10275 ( .A(n3469), .B(n3470), .C(n3471), .D(n3472), .Z(
        n3468) );
  HS65_LL_MX41X7 U10276 ( .D0(n193), .S0(n220), .D1(n209), .S1(n198), .D2(n219), .S2(n190), .D3(n203), .S3(n217), .Z(n3467) );
  HS65_LL_AOI212X4 U10277 ( .A(n221), .B(n3473), .C(n195), .D(n208), .E(n3474), 
        .Z(n3466) );
  HS65_LL_NOR4ABX2 U10278 ( .A(n3706), .B(n3707), .C(n3708), .D(n3709), .Z(
        n2976) );
  HS65_LL_NAND4ABX3 U10279 ( .A(n3710), .B(n3711), .C(n3712), .D(n3713), .Z(
        n3709) );
  HS65_LL_MX41X7 U10280 ( .D0(n636), .S0(n649), .D1(n658), .S1(n631), .D2(n651), .S2(n639), .D3(n625), .S3(n647), .Z(n3708) );
  HS65_LL_AOI212X4 U10281 ( .A(n650), .B(n3714), .C(n634), .D(n657), .E(n3715), 
        .Z(n3707) );
  HS65_LL_NOR4ABX2 U10282 ( .A(n8980), .B(n8981), .C(n8982), .D(n8983), .Z(
        n8642) );
  HS65_LL_NAND4ABX3 U10283 ( .A(n8209), .B(n7968), .C(n8286), .D(n8246), .Z(
        n8983) );
  HS65_LL_MX41X7 U10284 ( .D0(n363), .S0(n394), .D1(n378), .S1(n396), .D2(n390), .S2(n376), .D3(n395), .S3(n377), .Z(n8982) );
  HS65_LL_NOR4ABX2 U10285 ( .A(n8300), .B(n8098), .C(n8233), .D(n7984), .Z(
        n8980) );
  HS65_LL_NAND4ABX3 U10286 ( .A(n1786), .B(n1787), .C(n1788), .D(n1789), .Z(
        n1766) );
  HS65_LL_NAND4ABX3 U10287 ( .A(n1665), .B(n1541), .C(n1727), .D(n1686), .Z(
        n1787) );
  HS65_LL_NOR4ABX2 U10288 ( .A(n1618), .B(n1705), .C(n1648), .D(n1625), .Z(
        n1789) );
  HS65_LL_NOR4ABX2 U10289 ( .A(n1740), .B(n1563), .C(n1673), .D(n1603), .Z(
        n1788) );
  HS65_LL_NAND4ABX3 U10290 ( .A(n2162), .B(n2163), .C(n2164), .D(n2165), .Z(
        n2142) );
  HS65_LL_NAND4ABX3 U10291 ( .A(n2041), .B(n1917), .C(n2103), .D(n2062), .Z(
        n2163) );
  HS65_LL_NOR4ABX2 U10292 ( .A(n1994), .B(n2081), .C(n2024), .D(n2001), .Z(
        n2165) );
  HS65_LL_NOR4ABX2 U10293 ( .A(n2116), .B(n1939), .C(n2049), .D(n1979), .Z(
        n2164) );
  HS65_LL_NAND4ABX3 U10294 ( .A(n1410), .B(n1411), .C(n1412), .D(n1413), .Z(
        n1390) );
  HS65_LL_NAND4ABX3 U10295 ( .A(n1289), .B(n1165), .C(n1351), .D(n1310), .Z(
        n1411) );
  HS65_LL_NOR4ABX2 U10296 ( .A(n1242), .B(n1329), .C(n1272), .D(n1249), .Z(
        n1413) );
  HS65_LL_NOR4ABX2 U10297 ( .A(n1364), .B(n1187), .C(n1297), .D(n1227), .Z(
        n1412) );
  HS65_LL_NAND4ABX3 U10298 ( .A(n2538), .B(n2539), .C(n2540), .D(n2541), .Z(
        n2518) );
  HS65_LL_NAND4ABX3 U10299 ( .A(n2417), .B(n2293), .C(n2479), .D(n2438), .Z(
        n2539) );
  HS65_LL_NOR4ABX2 U10300 ( .A(n2370), .B(n2457), .C(n2400), .D(n2377), .Z(
        n2541) );
  HS65_LL_NOR4ABX2 U10301 ( .A(n2492), .B(n2315), .C(n2425), .D(n2355), .Z(
        n2540) );
  HS65_LL_NOR4ABX2 U10302 ( .A(n4133), .B(n4134), .C(n4135), .D(n4136), .Z(
        n4081) );
  HS65_LL_OR4X4 U10303 ( .A(n3277), .B(n3028), .C(n3234), .D(n3250), .Z(n4136)
         );
  HS65_LL_NAND4ABX3 U10304 ( .A(n3612), .B(n3650), .C(n3628), .D(n3596), .Z(
        n4135) );
  HS65_LL_AOI222X2 U10305 ( .A(n145), .B(n169), .C(n158), .D(n166), .E(n156), 
        .F(n174), .Z(n4133) );
  HS65_LL_NOR4ABX2 U10306 ( .A(n9068), .B(n9069), .C(n9070), .D(n9071), .Z(
        n7717) );
  HS65_LL_NAND4ABX3 U10307 ( .A(n8463), .B(n8826), .C(n8766), .D(n8450), .Z(
        n9071) );
  HS65_LL_NAND4ABX3 U10308 ( .A(n8792), .B(n8838), .C(n8171), .D(n8780), .Z(
        n9070) );
  HS65_LL_AOI222X2 U10309 ( .A(n102), .B(n127), .C(n134), .D(n113), .E(n112), 
        .F(n130), .Z(n9068) );
  HS65_LL_NOR4ABX2 U10310 ( .A(n9010), .B(n9011), .C(n9012), .D(n9013), .Z(
        n7679) );
  HS65_LL_NAND4ABX3 U10311 ( .A(n8411), .B(n8736), .C(n8676), .D(n8398), .Z(
        n9013) );
  HS65_LL_NAND4ABX3 U10312 ( .A(n8702), .B(n8748), .C(n8148), .D(n8690), .Z(
        n9012) );
  HS65_LL_AOI222X2 U10313 ( .A(n582), .B(n607), .C(n614), .D(n593), .E(n592), 
        .F(n610), .Z(n9010) );
  HS65_LL_NOR4ABX2 U10314 ( .A(n4010), .B(n4011), .C(n4012), .D(n4013), .Z(
        n3947) );
  HS65_LL_NAND4ABX3 U10315 ( .A(n3724), .B(n3137), .C(n3701), .D(n3763), .Z(
        n4013) );
  HS65_LL_MX41X7 U10316 ( .D0(n640), .S0(n649), .D1(n631), .S1(n651), .D2(n658), .S2(n630), .D3(n652), .S3(n628), .Z(n4012) );
  HS65_LL_NOR4ABX2 U10317 ( .A(n3334), .B(n3741), .C(n3672), .D(n3346), .Z(
        n4011) );
  HS65_LL_NOR4ABX2 U10318 ( .A(n8228), .B(n8229), .C(n8230), .D(n8231), .Z(
        n7862) );
  HS65_LL_NAND4ABX3 U10319 ( .A(n8232), .B(n8233), .C(n8234), .D(n8235), .Z(
        n8231) );
  HS65_LL_MX41X7 U10320 ( .D0(n369), .S0(n394), .D1(n390), .S1(n378), .D2(n396), .S2(n365), .D3(n372), .S3(n385), .Z(n8230) );
  HS65_LL_AOI212X4 U10321 ( .A(n393), .B(n8236), .C(n368), .D(n388), .E(n8237), 
        .Z(n8229) );
  HS65_LL_NOR4ABX2 U10322 ( .A(n4033), .B(n4034), .C(n4035), .D(n4036), .Z(
        n3967) );
  HS65_LL_NAND4ABX3 U10323 ( .A(n3815), .B(n3200), .C(n3878), .D(n3838), .Z(
        n4036) );
  HS65_LL_MX41X7 U10324 ( .D0(n422), .S0(n440), .D1(n413), .S1(n442), .D2(n427), .S2(n412), .D3(n443), .S3(n409), .Z(n4035) );
  HS65_LL_NOR4ABX2 U10325 ( .A(n3804), .B(n3177), .C(n3826), .D(n3374), .Z(
        n4033) );
  HS65_LL_NAND3X5 U10326 ( .A(n2531), .B(n2532), .C(n2533), .Z(n2253) );
  HS65_LL_NOR3AX2 U10327 ( .A(n2358), .B(n2485), .C(n2463), .Z(n2532) );
  HS65_LL_NOR3X4 U10328 ( .A(n2403), .B(n2537), .C(n2443), .Z(n2531) );
  HS65_LL_AOI212X4 U10329 ( .A(n885), .B(n914), .C(n904), .D(n880), .E(n2534), 
        .Z(n2533) );
  HS65_LL_NAND4ABX3 U10330 ( .A(n4192), .B(n4193), .C(n4194), .D(n4195), .Z(
        n3921) );
  HS65_LL_NAND4ABX3 U10331 ( .A(n3458), .B(n2935), .C(n3524), .D(n3483), .Z(
        n4193) );
  HS65_LL_MX41X7 U10332 ( .D0(n189), .S0(n220), .D1(n198), .S1(n219), .D2(n209), .S2(n199), .D3(n218), .S3(n196), .Z(n4192) );
  HS65_LL_NOR4ABX2 U10333 ( .A(n3106), .B(n3501), .C(n3429), .D(n3119), .Z(
        n4195) );
  HS65_LL_NOR4ABX2 U10334 ( .A(n2212), .B(n2213), .C(n2214), .D(n2215), .Z(
        n2141) );
  HS65_LL_NAND4ABX3 U10335 ( .A(n2000), .B(n2048), .C(n2117), .D(n1978), .Z(
        n2215) );
  HS65_LL_NAND4ABX3 U10336 ( .A(n1941), .B(n2064), .C(n2043), .D(n2080), .Z(
        n2214) );
  HS65_LL_AOI222X2 U10337 ( .A(n766), .B(n780), .C(n762), .D(n792), .E(n778), 
        .F(n769), .Z(n2212) );
  HS65_LL_NOR4ABX2 U10338 ( .A(n1460), .B(n1461), .C(n1462), .D(n1463), .Z(
        n1389) );
  HS65_LL_NAND4ABX3 U10339 ( .A(n1248), .B(n1296), .C(n1365), .D(n1226), .Z(
        n1463) );
  HS65_LL_NAND4ABX3 U10340 ( .A(n1189), .B(n1312), .C(n1291), .D(n1328), .Z(
        n1462) );
  HS65_LL_AOI222X2 U10341 ( .A(n848), .B(n862), .C(n844), .D(n874), .E(n860), 
        .F(n851), .Z(n1460) );
  HS65_LL_NOR4ABX2 U10342 ( .A(n1836), .B(n1837), .C(n1838), .D(n1839), .Z(
        n1765) );
  HS65_LL_NAND4ABX3 U10343 ( .A(n1624), .B(n1672), .C(n1741), .D(n1602), .Z(
        n1839) );
  HS65_LL_AOI222X2 U10344 ( .A(n807), .B(n821), .C(n803), .D(n833), .E(n819), 
        .F(n810), .Z(n1836) );
  HS65_LL_NAND4ABX3 U10345 ( .A(n1565), .B(n1688), .C(n1667), .D(n1704), .Z(
        n1838) );
  HS65_LL_NOR4ABX2 U10346 ( .A(n2588), .B(n2589), .C(n2590), .D(n2591), .Z(
        n2517) );
  HS65_LL_NAND4ABX3 U10347 ( .A(n2376), .B(n2424), .C(n2493), .D(n2354), .Z(
        n2591) );
  HS65_LL_NAND4ABX3 U10348 ( .A(n2317), .B(n2440), .C(n2419), .D(n2456), .Z(
        n2590) );
  HS65_LL_AOI222X2 U10349 ( .A(n889), .B(n903), .C(n885), .D(n915), .E(n901), 
        .F(n892), .Z(n2588) );
  HS65_LL_NOR4ABX2 U10350 ( .A(n4196), .B(n4197), .C(n4198), .D(n4199), .Z(
        n4050) );
  HS65_LL_NAND4ABX3 U10351 ( .A(n3118), .B(n3469), .C(n3448), .D(n3088), .Z(
        n4199) );
  HS65_LL_NAND4ABX3 U10352 ( .A(n2952), .B(n3485), .C(n3460), .D(n3500), .Z(
        n4198) );
  HS65_LL_AOI222X2 U10353 ( .A(n216), .B(n190), .C(n221), .D(n203), .E(n201), 
        .F(n212), .Z(n4196) );
  HS65_LL_NAND2X7 U10354 ( .A(n392), .B(n375), .Z(n8227) );
  HS65_LL_NAND4ABX3 U10355 ( .A(n3736), .B(n3737), .C(n3738), .D(n3739), .Z(
        n3313) );
  HS65_LL_NOR3AX2 U10356 ( .A(n3743), .B(n3744), .C(n3745), .Z(n3738) );
  HS65_LL_NAND4ABX3 U10357 ( .A(n3751), .B(n3752), .C(n3753), .D(n3754), .Z(
        n3736) );
  HS65_LL_NOR4ABX2 U10358 ( .A(n3740), .B(n3741), .C(n3742), .D(n2891), .Z(
        n3739) );
  HS65_LL_NAND4ABX3 U10359 ( .A(n8258), .B(n8259), .C(n8260), .D(n8261), .Z(
        n8092) );
  HS65_LL_NOR4ABX2 U10360 ( .A(n8266), .B(n8267), .C(n8268), .D(n8269), .Z(
        n8260) );
  HS65_LL_OR4X4 U10361 ( .A(n8274), .B(n8275), .C(n8276), .D(n7746), .Z(n8258)
         );
  HS65_LL_NOR4ABX2 U10362 ( .A(n8262), .B(n8263), .C(n8264), .D(n8265), .Z(
        n8261) );
  HS65_LL_NOR4ABX2 U10363 ( .A(n5625), .B(n5626), .C(n5627), .D(n5628), .Z(
        n5551) );
  HS65_LL_NAND4ABX3 U10364 ( .A(n5432), .B(n4797), .C(n5411), .D(n5386), .Z(
        n5628) );
  HS65_LL_MX41X7 U10365 ( .D0(n464), .S0(n473), .D1(n451), .S1(n476), .D2(n485), .S2(n452), .D3(n475), .S3(n449), .Z(n5627) );
  HS65_LL_NOR4ABX2 U10366 ( .A(n5443), .B(n4977), .C(n5366), .D(n4782), .Z(
        n5625) );
  HS65_LL_NOR4ABX2 U10367 ( .A(n5600), .B(n5601), .C(n5602), .D(n5603), .Z(
        n5529) );
  HS65_LL_NAND4ABX3 U10368 ( .A(n5317), .B(n4736), .C(n5296), .D(n5271), .Z(
        n5603) );
  HS65_LL_MX41X7 U10369 ( .D0(n247), .S0(n256), .D1(n234), .S1(n259), .D2(n268), .S2(n235), .D3(n258), .S3(n232), .Z(n5602) );
  HS65_LL_NOR4ABX2 U10370 ( .A(n5328), .B(n4924), .C(n5251), .D(n4755), .Z(
        n5600) );
  HS65_LL_NOR4ABX2 U10371 ( .A(n7217), .B(n7218), .C(n7219), .D(n7220), .Z(
        n7143) );
  HS65_LL_NAND4ABX3 U10372 ( .A(n7024), .B(n6390), .C(n7003), .D(n6978), .Z(
        n7220) );
  HS65_LL_MX41X7 U10373 ( .D0(n289), .S0(n298), .D1(n276), .S1(n301), .D2(n310), .S2(n277), .D3(n300), .S3(n274), .Z(n7219) );
  HS65_LL_NOR4ABX2 U10374 ( .A(n7035), .B(n6570), .C(n6958), .D(n6375), .Z(
        n7217) );
  HS65_LL_NOR4ABX2 U10375 ( .A(n5729), .B(n5730), .C(n5731), .D(n5732), .Z(
        n5504) );
  HS65_LL_NAND4ABX3 U10376 ( .A(n5079), .B(n4574), .C(n5058), .D(n5032), .Z(
        n5732) );
  HS65_LL_MX41X7 U10377 ( .D0(n10), .S0(n31), .D1(n24), .S1(n30), .D2(n39), 
        .S2(n25), .D3(n29), .S3(n22), .Z(n5731) );
  HS65_LL_NOR4ABX2 U10378 ( .A(n5106), .B(n4713), .C(n5011), .D(n4559), .Z(
        n5729) );
  HS65_LL_NOR4ABX2 U10379 ( .A(n5791), .B(n5792), .C(n5793), .D(n5794), .Z(
        n5568) );
  HS65_LL_NAND4ABX3 U10380 ( .A(n5201), .B(n4651), .C(n5180), .D(n5154), .Z(
        n5794) );
  HS65_LL_MX41X7 U10381 ( .D0(n666), .S0(n686), .D1(n679), .S1(n685), .D2(n694), .S2(n680), .D3(n684), .S3(n677), .Z(n5793) );
  HS65_LL_NOR4ABX2 U10382 ( .A(n5212), .B(n4851), .C(n5133), .D(n4636), .Z(
        n5791) );
  HS65_LL_NOR4ABX2 U10383 ( .A(n7383), .B(n7384), .C(n7385), .D(n7386), .Z(
        n7160) );
  HS65_LL_NAND4ABX3 U10384 ( .A(n6793), .B(n6244), .C(n6772), .D(n6746), .Z(
        n7386) );
  HS65_LL_MX41X7 U10385 ( .D0(n490), .S0(n510), .D1(n503), .S1(n509), .D2(n518), .S2(n504), .D3(n508), .S3(n501), .Z(n7385) );
  HS65_LL_NOR4ABX2 U10386 ( .A(n6804), .B(n6444), .C(n6725), .D(n6229), .Z(
        n7383) );
  HS65_LL_NOR4ABX2 U10387 ( .A(n7321), .B(n7322), .C(n7323), .D(n7324), .Z(
        n7096) );
  HS65_LL_NAND4ABX3 U10388 ( .A(n6672), .B(n6167), .C(n6651), .D(n6625), .Z(
        n7324) );
  HS65_LL_MX41X7 U10389 ( .D0(n532), .S0(n553), .D1(n546), .S1(n552), .D2(n561), .S2(n547), .D3(n551), .S3(n544), .Z(n7323) );
  HS65_LL_NOR4ABX2 U10390 ( .A(n6699), .B(n6306), .C(n6604), .D(n6152), .Z(
        n7321) );
  HS65_LL_NOR4ABX2 U10391 ( .A(n7192), .B(n7193), .C(n7194), .D(n7195), .Z(
        n7121) );
  HS65_LL_NAND4ABX3 U10392 ( .A(n6909), .B(n6351), .C(n6888), .D(n6863), .Z(
        n7195) );
  HS65_LL_MX41X7 U10393 ( .D0(n68), .S0(n74), .D1(n63), .S1(n77), .D2(n82), 
        .S2(n66), .D3(n73), .S3(n65), .Z(n7194) );
  HS65_LL_NOR4ABX2 U10394 ( .A(n6920), .B(n6517), .C(n6843), .D(n6336), .Z(
        n7192) );
  HS65_LL_NAND4ABX3 U10395 ( .A(n2452), .B(n2453), .C(n2454), .D(n2455), .Z(
        n2348) );
  HS65_LL_NOR3AX2 U10396 ( .A(n2459), .B(n2460), .C(n2461), .Z(n2454) );
  HS65_LL_NAND4ABX3 U10397 ( .A(n2463), .B(n2464), .C(n2465), .D(n2466), .Z(
        n2453) );
  HS65_LL_NOR4ABX2 U10398 ( .A(n2456), .B(n2457), .C(n2458), .D(n2247), .Z(
        n2455) );
  HS65_LL_NAND4ABX3 U10399 ( .A(n1324), .B(n1325), .C(n1326), .D(n1327), .Z(
        n1220) );
  HS65_LL_NAND4ABX3 U10400 ( .A(n1335), .B(n1336), .C(n1337), .D(n1338), .Z(
        n1325) );
  HS65_LL_NOR3AX2 U10401 ( .A(n1331), .B(n1332), .C(n1333), .Z(n1326) );
  HS65_LL_NOR4ABX2 U10402 ( .A(n1328), .B(n1329), .C(n1330), .D(n1119), .Z(
        n1327) );
  HS65_LL_NAND4ABX3 U10403 ( .A(n2076), .B(n2077), .C(n2078), .D(n2079), .Z(
        n1972) );
  HS65_LL_NAND4ABX3 U10404 ( .A(n2087), .B(n2088), .C(n2089), .D(n2090), .Z(
        n2077) );
  HS65_LL_NOR3AX2 U10405 ( .A(n2083), .B(n2084), .C(n2085), .Z(n2078) );
  HS65_LL_NOR4ABX2 U10406 ( .A(n2080), .B(n2081), .C(n2082), .D(n1871), .Z(
        n2079) );
  HS65_LL_NAND4ABX3 U10407 ( .A(n1700), .B(n1701), .C(n1702), .D(n1703), .Z(
        n1596) );
  HS65_LL_NOR3AX2 U10408 ( .A(n1707), .B(n1708), .C(n1709), .Z(n1702) );
  HS65_LL_NOR4ABX2 U10409 ( .A(n1704), .B(n1705), .C(n1706), .D(n1495), .Z(
        n1703) );
  HS65_LL_NAND4ABX3 U10410 ( .A(n1711), .B(n1712), .C(n1713), .D(n1714), .Z(
        n1701) );
  HS65_LL_NAND4ABX3 U10411 ( .A(n3851), .B(n3852), .C(n3853), .D(n3854), .Z(
        n3367) );
  HS65_LL_NOR3AX2 U10412 ( .A(n3858), .B(n3859), .C(n3860), .Z(n3853) );
  HS65_LL_NOR4ABX2 U10413 ( .A(n3855), .B(n3856), .C(n3857), .D(n2839), .Z(
        n3854) );
  HS65_LL_NAND4ABX3 U10414 ( .A(n3866), .B(n3867), .C(n3868), .D(n3869), .Z(
        n3851) );
  HS65_LL_NAND4ABX3 U10415 ( .A(n3496), .B(n3497), .C(n3498), .D(n3499), .Z(
        n3082) );
  HS65_LL_NOR3AX2 U10416 ( .A(n3504), .B(n3505), .C(n3506), .Z(n3498) );
  HS65_LL_NAND4ABX3 U10417 ( .A(n3508), .B(n3509), .C(n3510), .D(n3511), .Z(
        n3497) );
  HS65_LL_NOR4ABX2 U10418 ( .A(n3500), .B(n3501), .C(n3502), .D(n3503), .Z(
        n3499) );
  HS65_LL_NOR4ABX2 U10419 ( .A(n8912), .B(n8913), .C(n8914), .D(n8915), .Z(
        n8855) );
  HS65_LL_NAND4ABX3 U10420 ( .A(n8512), .B(n8589), .C(n8037), .D(n8548), .Z(
        n8915) );
  HS65_LL_MX41X7 U10421 ( .D0(n320), .S0(n354), .D1(n330), .S1(n356), .D2(n342), .S2(n328), .D3(n353), .S3(n329), .Z(n8914) );
  HS65_LL_NOR4ABX2 U10422 ( .A(n8525), .B(n8331), .C(n8535), .D(n8052), .Z(
        n8912) );
  HS65_LL_NOR4ABX2 U10423 ( .A(n2420), .B(n2421), .C(n2422), .D(n2423), .Z(
        n2266) );
  HS65_LL_MX41X7 U10424 ( .D0(n904), .S0(n890), .D1(n888), .S1(n907), .D2(n895), .S2(n903), .D3(n915), .S3(n2428), .Z(n2422) );
  HS65_LL_NAND4ABX3 U10425 ( .A(n2424), .B(n2425), .C(n2426), .D(n2427), .Z(
        n2423) );
  HS65_LL_AOI212X4 U10426 ( .A(n885), .B(n2429), .C(n910), .D(n887), .E(n2430), 
        .Z(n2421) );
  HS65_LL_NOR4ABX2 U10427 ( .A(n1292), .B(n1293), .C(n1294), .D(n1295), .Z(
        n1138) );
  HS65_LL_MX41X7 U10428 ( .D0(n863), .S0(n849), .D1(n847), .S1(n866), .D2(n854), .S2(n862), .D3(n874), .S3(n1300), .Z(n1294) );
  HS65_LL_NAND4ABX3 U10429 ( .A(n1296), .B(n1297), .C(n1298), .D(n1299), .Z(
        n1295) );
  HS65_LL_AOI212X4 U10430 ( .A(n844), .B(n1301), .C(n869), .D(n846), .E(n1302), 
        .Z(n1293) );
  HS65_LL_NOR4ABX2 U10431 ( .A(n1668), .B(n1669), .C(n1670), .D(n1671), .Z(
        n1514) );
  HS65_LL_MX41X7 U10432 ( .D0(n822), .S0(n808), .D1(n806), .S1(n825), .D2(n813), .S2(n821), .D3(n833), .S3(n1676), .Z(n1670) );
  HS65_LL_NAND4ABX3 U10433 ( .A(n1672), .B(n1673), .C(n1674), .D(n1675), .Z(
        n1671) );
  HS65_LL_AOI212X4 U10434 ( .A(n803), .B(n1677), .C(n828), .D(n805), .E(n1678), 
        .Z(n1669) );
  HS65_LL_NOR4ABX2 U10435 ( .A(n2044), .B(n2045), .C(n2046), .D(n2047), .Z(
        n1890) );
  HS65_LL_MX41X7 U10436 ( .D0(n781), .S0(n767), .D1(n765), .S1(n784), .D2(n772), .S2(n780), .D3(n792), .S3(n2052), .Z(n2046) );
  HS65_LL_NAND4ABX3 U10437 ( .A(n2048), .B(n2049), .C(n2050), .D(n2051), .Z(
        n2047) );
  HS65_LL_AOI212X4 U10438 ( .A(n762), .B(n2053), .C(n787), .D(n764), .E(n2054), 
        .Z(n2045) );
  HS65_LL_NAND2X7 U10439 ( .A(n37), .B(n14), .Z(n4721) );
  HS65_LL_NAND2X7 U10440 ( .A(n559), .B(n536), .Z(n6314) );
  HS65_LL_NAND4ABX3 U10441 ( .A(n8691), .B(n8692), .C(n8693), .D(n8694), .Z(
        n8386) );
  HS65_LL_NOR4ABX2 U10442 ( .A(n7692), .B(n7625), .C(n7798), .D(n8695), .Z(
        n8694) );
  HS65_LL_NOR4ABX2 U10443 ( .A(n8696), .B(n8697), .C(n8698), .D(n7826), .Z(
        n8693) );
  HS65_LL_NAND4ABX3 U10444 ( .A(n8702), .B(n8703), .C(n7815), .D(n7670), .Z(
        n8691) );
  HS65_LL_NAND4ABX3 U10445 ( .A(n8781), .B(n8782), .C(n8783), .D(n8784), .Z(
        n8438) );
  HS65_LL_NOR4ABX2 U10446 ( .A(n7730), .B(n7665), .C(n7897), .D(n8785), .Z(
        n8784) );
  HS65_LL_NOR4ABX2 U10447 ( .A(n8786), .B(n8787), .C(n8788), .D(n7924), .Z(
        n8783) );
  HS65_LL_NAND4ABX3 U10448 ( .A(n8792), .B(n8793), .C(n7913), .D(n7708), .Z(
        n8781) );
  HS65_LL_NAND2X7 U10449 ( .A(n100), .B(n136), .Z(n8450) );
  HS65_LL_NAND2X7 U10450 ( .A(n152), .B(n178), .Z(n3544) );
  HS65_LL_NOR2X6 U10451 ( .A(n850), .B(n852), .Z(n1155) );
  HS65_LL_NAND4ABX3 U10452 ( .A(n2578), .B(n2579), .C(n2580), .D(n2581), .Z(
        n2508) );
  HS65_LL_NAND4ABX3 U10453 ( .A(n2392), .B(n2345), .C(n2584), .D(n2405), .Z(
        n2579) );
  HS65_LL_AOI222X2 U10454 ( .A(n896), .B(n903), .C(n907), .D(n880), .E(n888), 
        .F(n915), .Z(n2580) );
  HS65_LL_NOR4ABX2 U10455 ( .A(n2363), .B(n2475), .C(n2449), .D(n2468), .Z(
        n2581) );
  HS65_LL_NAND4ABX3 U10456 ( .A(n2202), .B(n2203), .C(n2204), .D(n2205), .Z(
        n2132) );
  HS65_LL_AOI222X2 U10457 ( .A(n773), .B(n780), .C(n784), .D(n757), .E(n765), 
        .F(n792), .Z(n2204) );
  HS65_LL_NAND4ABX3 U10458 ( .A(n2016), .B(n1969), .C(n2208), .D(n2029), .Z(
        n2203) );
  HS65_LL_NOR4ABX2 U10459 ( .A(n1987), .B(n2099), .C(n2073), .D(n2092), .Z(
        n2205) );
  HS65_LL_NAND4ABX3 U10460 ( .A(n1826), .B(n1827), .C(n1828), .D(n1829), .Z(
        n1756) );
  HS65_LL_AOI222X2 U10461 ( .A(n814), .B(n821), .C(n825), .D(n798), .E(n806), 
        .F(n833), .Z(n1828) );
  HS65_LL_NAND4ABX3 U10462 ( .A(n1640), .B(n1593), .C(n1832), .D(n1653), .Z(
        n1827) );
  HS65_LL_NOR4ABX2 U10463 ( .A(n1611), .B(n1723), .C(n1697), .D(n1716), .Z(
        n1829) );
  HS65_LL_NAND4ABX3 U10464 ( .A(n1450), .B(n1451), .C(n1452), .D(n1453), .Z(
        n1380) );
  HS65_LL_AOI222X2 U10465 ( .A(n855), .B(n862), .C(n866), .D(n839), .E(n847), 
        .F(n874), .Z(n1452) );
  HS65_LL_NAND4ABX3 U10466 ( .A(n1264), .B(n1217), .C(n1456), .D(n1277), .Z(
        n1451) );
  HS65_LL_NOR4ABX2 U10467 ( .A(n1235), .B(n1347), .C(n1321), .D(n1340), .Z(
        n1453) );
  HS65_LL_NAND4ABX3 U10468 ( .A(n2393), .B(n2394), .C(n2395), .D(n2396), .Z(
        n2347) );
  HS65_LL_NOR4ABX2 U10469 ( .A(n2401), .B(n2402), .C(n2403), .D(n2404), .Z(
        n2395) );
  HS65_LL_NOR4ABX2 U10470 ( .A(n2397), .B(n2398), .C(n2399), .D(n2400), .Z(
        n2396) );
  HS65_LL_NAND3X5 U10471 ( .A(n2405), .B(n2406), .C(n2407), .Z(n2393) );
  HS65_LL_NAND2X7 U10472 ( .A(n238), .B(n253), .Z(n4932) );
  HS65_LL_NAND2X7 U10473 ( .A(n455), .B(n470), .Z(n4985) );
  HS65_LL_NAND2X7 U10474 ( .A(n280), .B(n295), .Z(n6578) );
  HS65_LL_NAND2X7 U10475 ( .A(n60), .B(n88), .Z(n6525) );
  HS65_LL_NAND4ABX3 U10476 ( .A(n2017), .B(n2018), .C(n2019), .D(n2020), .Z(
        n1971) );
  HS65_LL_NOR4ABX2 U10477 ( .A(n2025), .B(n2026), .C(n2027), .D(n2028), .Z(
        n2019) );
  HS65_LL_NOR4ABX2 U10478 ( .A(n2021), .B(n2022), .C(n2023), .D(n2024), .Z(
        n2020) );
  HS65_LL_NAND3X5 U10479 ( .A(n2029), .B(n2030), .C(n2031), .Z(n2017) );
  HS65_LL_NAND4ABX3 U10480 ( .A(n1265), .B(n1266), .C(n1267), .D(n1268), .Z(
        n1219) );
  HS65_LL_NOR4ABX2 U10481 ( .A(n1273), .B(n1274), .C(n1275), .D(n1276), .Z(
        n1267) );
  HS65_LL_NOR4ABX2 U10482 ( .A(n1269), .B(n1270), .C(n1271), .D(n1272), .Z(
        n1268) );
  HS65_LL_NAND3X5 U10483 ( .A(n1277), .B(n1278), .C(n1279), .Z(n1265) );
  HS65_LL_NAND4ABX3 U10484 ( .A(n1641), .B(n1642), .C(n1643), .D(n1644), .Z(
        n1595) );
  HS65_LL_NOR4ABX2 U10485 ( .A(n1649), .B(n1650), .C(n1651), .D(n1652), .Z(
        n1643) );
  HS65_LL_NOR4ABX2 U10486 ( .A(n1645), .B(n1646), .C(n1647), .D(n1648), .Z(
        n1644) );
  HS65_LL_MX41X7 U10487 ( .D0(n822), .S0(n810), .D1(n819), .S1(n798), .D2(n799), .S2(n832), .D3(n800), .S3(n830), .Z(n1642) );
  HS65_LL_NAND4ABX3 U10488 ( .A(n3780), .B(n3781), .C(n3782), .D(n3783), .Z(
        n3366) );
  HS65_LL_NOR4ABX2 U10489 ( .A(n3788), .B(n3789), .C(n3790), .D(n3791), .Z(
        n3782) );
  HS65_LL_NOR4ABX2 U10490 ( .A(n3784), .B(n3785), .C(n3786), .D(n3787), .Z(
        n3783) );
  HS65_LL_NAND3AX6 U10491 ( .A(n3792), .B(n3793), .C(n3794), .Z(n3780) );
  HS65_LL_NAND4ABX3 U10492 ( .A(n3665), .B(n3666), .C(n3667), .D(n3668), .Z(
        n3312) );
  HS65_LL_NOR4ABX2 U10493 ( .A(n3673), .B(n3674), .C(n3675), .D(n3676), .Z(
        n3667) );
  HS65_LL_NAND3AX6 U10494 ( .A(n3677), .B(n3678), .C(n3679), .Z(n3665) );
  HS65_LL_NOR4ABX2 U10495 ( .A(n3669), .B(n3670), .C(n3671), .D(n3672), .Z(
        n3668) );
  HS65_LL_NAND2X7 U10496 ( .A(n400), .B(n374), .Z(n7970) );
  HS65_LL_NOR2X6 U10497 ( .A(n763), .B(n758), .Z(n1901) );
  HS65_LL_NAND2X7 U10498 ( .A(n770), .B(n785), .Z(n2029) );
  HS65_LL_NAND2X7 U10499 ( .A(n811), .B(n826), .Z(n1653) );
  HS65_LL_NAND2X7 U10500 ( .A(n893), .B(n908), .Z(n2405) );
  HS65_LL_NAND2X7 U10501 ( .A(n852), .B(n867), .Z(n1277) );
  HS65_LL_NAND2X7 U10502 ( .A(n324), .B(n351), .Z(n8548) );
  HS65_LL_NOR2X6 U10503 ( .A(n886), .B(n881), .Z(n2277) );
  HS65_LL_NOR2X6 U10504 ( .A(n845), .B(n840), .Z(n1149) );
  HS65_LL_NAND2X7 U10505 ( .A(n327), .B(n355), .Z(n8601) );
  HS65_LL_NAND2X7 U10506 ( .A(n98), .B(n127), .Z(n7913) );
  HS65_LL_NAND2X7 U10507 ( .A(n578), .B(n607), .Z(n7815) );
  HS65_LL_NAND2X7 U10508 ( .A(n328), .B(n349), .Z(n8354) );
  HS65_LL_NAND2X7 U10509 ( .A(n454), .B(n485), .Z(n5411) );
  HS65_LL_NAND2X7 U10510 ( .A(n237), .B(n268), .Z(n5296) );
  HS65_LL_NAND2X7 U10511 ( .A(n279), .B(n310), .Z(n7003) );
  HS65_LL_NAND2X7 U10512 ( .A(n58), .B(n82), .Z(n6888) );
  HS65_LL_NAND2X7 U10513 ( .A(n914), .B(n890), .Z(n2493) );
  HS65_LL_NAND2X7 U10514 ( .A(n791), .B(n767), .Z(n2117) );
  HS65_LL_NAND2X7 U10515 ( .A(n873), .B(n849), .Z(n1365) );
  HS65_LL_NAND2X7 U10516 ( .A(n906), .B(n889), .Z(n2406) );
  HS65_LL_NAND2X7 U10517 ( .A(n832), .B(n808), .Z(n1741) );
  HS65_LL_NAND2X7 U10518 ( .A(n65), .B(n84), .Z(n6924) );
  HS65_LL_NAND2X7 U10519 ( .A(n232), .B(n262), .Z(n5332) );
  HS65_LL_NAND2X7 U10520 ( .A(n449), .B(n479), .Z(n5447) );
  HS65_LL_NAND2X7 U10521 ( .A(n274), .B(n304), .Z(n7039) );
  HS65_LL_NAND2X7 U10522 ( .A(n501), .B(n515), .Z(n6808) );
  HS65_LL_NAND2X7 U10523 ( .A(n417), .B(n440), .Z(n3805) );
  HS65_LL_NAND2X7 U10524 ( .A(n194), .B(n220), .Z(n3448) );
  HS65_LL_NAND2X7 U10525 ( .A(n865), .B(n848), .Z(n1278) );
  HS65_LL_NAND2X7 U10526 ( .A(n783), .B(n766), .Z(n2030) );
  HS65_LL_NAND2X7 U10527 ( .A(n824), .B(n807), .Z(n1654) );
  HS65_LL_NAND2X7 U10528 ( .A(n786), .B(n763), .Z(n2043) );
  HS65_LL_NAND2X7 U10529 ( .A(n868), .B(n845), .Z(n1291) );
  HS65_LL_NAND2X7 U10530 ( .A(n659), .B(n635), .Z(n3750) );
  HS65_LL_NAND2X7 U10531 ( .A(n904), .B(n889), .Z(n2465) );
  HS65_LL_NAND2X7 U10532 ( .A(n635), .B(n649), .Z(n3690) );
  HS65_LL_NAND2X7 U10533 ( .A(n909), .B(n886), .Z(n2419) );
  HS65_LL_NAND2X7 U10534 ( .A(n863), .B(n848), .Z(n1337) );
  HS65_LL_NAND2X7 U10535 ( .A(n781), .B(n766), .Z(n2089) );
  HS65_LL_NAND2X7 U10536 ( .A(n901), .B(n889), .Z(n2379) );
  HS65_LL_NAND2X7 U10537 ( .A(n811), .B(n824), .Z(n1617) );
  HS65_LL_NAND2X7 U10538 ( .A(n827), .B(n804), .Z(n1667) );
  HS65_LL_NAND2X7 U10539 ( .A(n822), .B(n807), .Z(n1713) );
  HS65_LL_NAND2X7 U10540 ( .A(n860), .B(n848), .Z(n1251) );
  HS65_LL_NAND2X7 U10541 ( .A(n778), .B(n766), .Z(n2003) );
  HS65_LL_NAND2X7 U10542 ( .A(n893), .B(n906), .Z(n2369) );
  HS65_LL_NAND2X7 U10543 ( .A(n770), .B(n783), .Z(n1993) );
  HS65_LL_NAND2X7 U10544 ( .A(n852), .B(n865), .Z(n1241) );
  HS65_LL_NAND2X7 U10545 ( .A(n819), .B(n807), .Z(n1627) );
  HS65_LL_NAND2X7 U10546 ( .A(n420), .B(n438), .Z(n3817) );
  HS65_LL_NOR4ABX2 U10547 ( .A(n3893), .B(n3918), .C(n3919), .D(n3920), .Z(
        n3917) );
  HS65_LL_AOI212X4 U10548 ( .A(n189), .B(n216), .C(n211), .D(n188), .E(n3921), 
        .Z(n3918) );
  HS65_LL_NOR4ABX2 U10549 ( .A(n1381), .B(n1401), .C(n1125), .D(n1402), .Z(
        n1400) );
  HS65_LL_AOI212X4 U10550 ( .A(n875), .B(n848), .C(n842), .D(n868), .E(n1390), 
        .Z(n1401) );
  HS65_LL_NOR4ABX2 U10551 ( .A(n2133), .B(n2153), .C(n1877), .D(n2154), .Z(
        n2152) );
  HS65_LL_AOI212X4 U10552 ( .A(n793), .B(n766), .C(n760), .D(n786), .E(n2142), 
        .Z(n2153) );
  HS65_LL_NOR4ABX2 U10553 ( .A(n1757), .B(n1777), .C(n1501), .D(n1778), .Z(
        n1776) );
  HS65_LL_AOI212X4 U10554 ( .A(n834), .B(n807), .C(n801), .D(n827), .E(n1766), 
        .Z(n1777) );
  HS65_LL_NOR4ABX2 U10555 ( .A(n2509), .B(n2529), .C(n2253), .D(n2530), .Z(
        n2528) );
  HS65_LL_AOI212X4 U10556 ( .A(n916), .B(n889), .C(n883), .D(n909), .E(n2518), 
        .Z(n2529) );
  HS65_LL_NAND2X7 U10557 ( .A(n193), .B(n216), .Z(n3510) );
  HS65_LL_NAND2X7 U10558 ( .A(n188), .B(n214), .Z(n3460) );
  HS65_LL_NAND2X7 U10559 ( .A(n460), .B(n473), .Z(n5442) );
  HS65_LL_NAND2X7 U10560 ( .A(n285), .B(n298), .Z(n7034) );
  HS65_LL_NOR4ABX2 U10561 ( .A(n5543), .B(n5544), .C(n5545), .D(n4511), .Z(
        n5542) );
  HS65_LL_AOI212X4 U10562 ( .A(n470), .B(n458), .C(n464), .D(n467), .E(n5557), 
        .Z(n5544) );
  HS65_LL_NOR4ABX2 U10563 ( .A(n5521), .B(n5522), .C(n5523), .D(n4450), .Z(
        n5520) );
  HS65_LL_AOI212X4 U10564 ( .A(n253), .B(n241), .C(n247), .D(n250), .E(n5535), 
        .Z(n5522) );
  HS65_LL_NOR4ABX2 U10565 ( .A(n7135), .B(n7136), .C(n7137), .D(n6104), .Z(
        n7134) );
  HS65_LL_AOI212X4 U10566 ( .A(n295), .B(n283), .C(n289), .D(n292), .E(n7149), 
        .Z(n7136) );
  HS65_LL_NOR4ABX2 U10567 ( .A(n7113), .B(n7114), .C(n7115), .D(n6043), .Z(
        n7112) );
  HS65_LL_AOI212X4 U10568 ( .A(n88), .B(n57), .C(n68), .D(n91), .E(n7127), .Z(
        n7114) );
  HS65_LL_NAND2X7 U10569 ( .A(n24), .B(n37), .Z(n5109) );
  HS65_LL_NAND2X7 U10570 ( .A(n546), .B(n559), .Z(n6702) );
  HS65_LL_NOR4ABX2 U10571 ( .A(n4961), .B(n4939), .C(n4767), .D(n4602), .Z(
        n5353) );
  HS65_LL_NOR4ABX2 U10572 ( .A(n6554), .B(n6532), .C(n6360), .D(n6195), .Z(
        n6945) );
  HS65_LL_NAND2X7 U10573 ( .A(n348), .B(n325), .Z(n8536) );
  HS65_LL_NAND2X7 U10574 ( .A(n387), .B(n374), .Z(n8234) );
  HS65_LL_NAND2X7 U10575 ( .A(n354), .B(n334), .Z(n8524) );
  HS65_LL_NAND2X7 U10576 ( .A(n394), .B(n370), .Z(n8299) );
  HS65_LL_NOR4ABX2 U10577 ( .A(n7678), .B(n7679), .C(n7680), .D(n7629), .Z(
        n7668) );
  HS65_LL_NOR4ABX2 U10578 ( .A(n7716), .B(n7717), .C(n7718), .D(n7649), .Z(
        n7706) );
  HS65_LL_NAND2X7 U10579 ( .A(n418), .B(n436), .Z(n3864) );
  HS65_LL_NAND2X7 U10580 ( .A(n661), .B(n637), .Z(n3702) );
  HS65_LL_NOR4ABX2 U10581 ( .A(n5509), .B(n5644), .C(n5645), .D(n5475), .Z(
        n5640) );
  HS65_LL_NOR4ABX2 U10582 ( .A(n5592), .B(n5528), .C(n4451), .D(n5523), .Z(
        n5821) );
  HS65_LL_NOR4ABX2 U10583 ( .A(n5617), .B(n5550), .C(n4512), .D(n5545), .Z(
        n5880) );
  HS65_LL_NOR4ABX2 U10584 ( .A(n5573), .B(n5674), .C(n5675), .D(n5489), .Z(
        n5670) );
  HS65_LL_NOR4ABX2 U10585 ( .A(n7209), .B(n7142), .C(n6105), .D(n7137), .Z(
        n7472) );
  HS65_LL_NOR4ABX2 U10586 ( .A(n7165), .B(n7266), .C(n7267), .D(n7081), .Z(
        n7262) );
  HS65_LL_NAND2X7 U10587 ( .A(n362), .B(n384), .Z(n8108) );
  HS65_LL_NAND4ABX3 U10588 ( .A(n1619), .B(n1620), .C(n1621), .D(n1622), .Z(
        n1516) );
  HS65_LL_NOR3X4 U10589 ( .A(n1623), .B(n1624), .C(n1625), .Z(n1622) );
  HS65_LL_NAND3AX6 U10590 ( .A(n1626), .B(n1627), .C(n1628), .Z(n1620) );
  HS65_LL_AOI222X2 U10591 ( .A(n824), .B(n804), .C(n822), .D(n806), .E(n828), 
        .F(n809), .Z(n1621) );
  HS65_LL_NAND4ABX3 U10592 ( .A(n2371), .B(n2372), .C(n2373), .D(n2374), .Z(
        n2268) );
  HS65_LL_NOR3X4 U10593 ( .A(n2375), .B(n2376), .C(n2377), .Z(n2374) );
  HS65_LL_AOI222X2 U10594 ( .A(n906), .B(n886), .C(n904), .D(n888), .E(n910), 
        .F(n891), .Z(n2373) );
  HS65_LL_NAND3AX6 U10595 ( .A(n2378), .B(n2379), .C(n2380), .Z(n2372) );
  HS65_LL_NAND4ABX3 U10596 ( .A(n1243), .B(n1244), .C(n1245), .D(n1246), .Z(
        n1140) );
  HS65_LL_NOR3X4 U10597 ( .A(n1247), .B(n1248), .C(n1249), .Z(n1246) );
  HS65_LL_AOI222X2 U10598 ( .A(n865), .B(n845), .C(n863), .D(n847), .E(n869), 
        .F(n850), .Z(n1245) );
  HS65_LL_NAND3AX6 U10599 ( .A(n1250), .B(n1251), .C(n1252), .Z(n1244) );
  HS65_LL_NAND4ABX3 U10600 ( .A(n1995), .B(n1996), .C(n1997), .D(n1998), .Z(
        n1892) );
  HS65_LL_NOR3X4 U10601 ( .A(n1999), .B(n2000), .C(n2001), .Z(n1998) );
  HS65_LL_AOI222X2 U10602 ( .A(n783), .B(n763), .C(n781), .D(n765), .E(n787), 
        .F(n768), .Z(n1997) );
  HS65_LL_NAND3AX6 U10603 ( .A(n2002), .B(n2003), .C(n2004), .Z(n1996) );
  HS65_LL_NAND2X7 U10604 ( .A(n415), .B(n436), .Z(n3793) );
  HS65_LL_NOR3AX2 U10605 ( .A(n3896), .B(n4051), .C(n3919), .Z(n4166) );
  HS65_LL_NOR4ABX2 U10606 ( .A(n2906), .B(n2907), .C(n2908), .D(n2909), .Z(
        n2905) );
  HS65_LL_AO212X4 U10607 ( .A(n148), .B(n166), .C(n180), .D(n143), .E(n2910), 
        .Z(n2908) );
  HS65_LL_NAND2X7 U10608 ( .A(n280), .B(n298), .Z(n6541) );
  HS65_LL_NAND2X7 U10609 ( .A(n455), .B(n473), .Z(n4948) );
  HS65_LL_NOR2X6 U10610 ( .A(n602), .B(n614), .Z(n8742) );
  HS65_LL_NOR3AX2 U10611 ( .A(n2878), .B(n2879), .C(n2880), .Z(n2872) );
  HS65_LL_NOR4ABX2 U10612 ( .A(n7771), .B(n8855), .C(n8856), .D(n8857), .Z(
        n8854) );
  HS65_LL_MX41X7 U10613 ( .D0(n333), .S0(n341), .D1(n325), .S1(n352), .D2(n353), .S2(n330), .D3(n327), .S3(n348), .Z(n8856) );
  HS65_LL_NOR4ABX2 U10614 ( .A(n7753), .B(n8642), .C(n8643), .D(n8644), .Z(
        n8641) );
  HS65_LL_MX41X7 U10615 ( .D0(n367), .S0(n391), .D1(n374), .S1(n397), .D2(n395), .S2(n378), .D3(n375), .S3(n387), .Z(n8643) );
  HS65_LL_NOR3AX2 U10616 ( .A(n2986), .B(n3356), .C(n3171), .Z(n3352) );
  HS65_LL_NOR4ABX2 U10617 ( .A(n4095), .B(n4081), .C(n3988), .D(n4128), .Z(
        n4127) );
  HS65_LL_MX41X7 U10618 ( .D0(n147), .S0(n173), .D1(n168), .S1(n157), .D2(n163), .S2(n153), .D3(n152), .S3(n179), .Z(n4128) );
  HS65_LL_NAND2X7 U10619 ( .A(n21), .B(n31), .Z(n4665) );
  HS65_LL_NAND2X7 U10620 ( .A(n543), .B(n553), .Z(n6258) );
  HS65_LL_NAND3X5 U10621 ( .A(n8886), .B(n8887), .C(n8888), .Z(n8857) );
  HS65_LL_NOR4ABX2 U10622 ( .A(n8332), .B(n8514), .C(n8345), .D(n8360), .Z(
        n8887) );
  HS65_LL_NOR4ABX2 U10623 ( .A(n8537), .B(n8547), .C(n7954), .D(n8522), .Z(
        n8886) );
  HS65_LL_NOR4ABX2 U10624 ( .A(n8587), .B(n8053), .C(n8889), .D(n8890), .Z(
        n8888) );
  HS65_LL_NAND2X7 U10625 ( .A(n782), .B(n768), .Z(n2093) );
  HS65_LL_NAND2X7 U10626 ( .A(n864), .B(n850), .Z(n1341) );
  HS65_LL_NOR4ABX2 U10627 ( .A(n7678), .B(n7626), .C(n8999), .D(n7800), .Z(
        n8998) );
  HS65_LL_AO212X4 U10628 ( .A(n600), .B(n579), .C(n583), .D(n603), .E(n7697), 
        .Z(n8999) );
  HS65_LL_NOR4ABX2 U10629 ( .A(n7716), .B(n7646), .C(n9057), .D(n7899), .Z(
        n9056) );
  HS65_LL_AO212X4 U10630 ( .A(n120), .B(n99), .C(n103), .D(n123), .E(n7735), 
        .Z(n9057) );
  HS65_LL_NAND2X7 U10631 ( .A(n905), .B(n891), .Z(n2469) );
  HS65_LL_NAND2X7 U10632 ( .A(n842), .B(n864), .Z(n1290) );
  HS65_LL_NAND2X7 U10633 ( .A(n760), .B(n782), .Z(n2042) );
  HS65_LL_NAND2X7 U10634 ( .A(n801), .B(n823), .Z(n1666) );
  HS65_LL_NAND2X7 U10635 ( .A(n883), .B(n905), .Z(n2418) );
  HS65_LL_NAND2X7 U10636 ( .A(n823), .B(n809), .Z(n1717) );
  HS65_LL_NOR4ABX2 U10637 ( .A(n4317), .B(n3879), .C(n3387), .D(n3786), .Z(
        n4316) );
  HS65_LL_OAI21X3 U10638 ( .A(n418), .B(n419), .C(n442), .Z(n4317) );
  HS65_LL_NOR4ABX2 U10639 ( .A(n4258), .B(n3335), .C(n3766), .D(n3671), .Z(
        n4257) );
  HS65_LL_OAI21X3 U10640 ( .A(n636), .B(n637), .C(n651), .Z(n4258) );
  HS65_LL_NOR4ABX2 U10641 ( .A(n1206), .B(n1138), .C(n1170), .D(n1219), .Z(
        n1258) );
  HS65_LL_NOR4ABX2 U10642 ( .A(n1958), .B(n1890), .C(n1922), .D(n1971), .Z(
        n2010) );
  HS65_LL_NOR4ABX2 U10643 ( .A(n2334), .B(n2266), .C(n2298), .D(n2347), .Z(
        n2386) );
  HS65_LL_NOR4ABX2 U10644 ( .A(n1582), .B(n1514), .C(n1546), .D(n1595), .Z(
        n1634) );
  HS65_LL_NOR2X6 U10645 ( .A(n894), .B(n885), .Z(n2496) );
  HS65_LL_NOR2X6 U10646 ( .A(n771), .B(n762), .Z(n2120) );
  HS65_LL_NOR4ABX2 U10647 ( .A(n2265), .B(n2266), .C(n2267), .D(n2268), .Z(
        n2264) );
  HS65_LL_AO212X4 U10648 ( .A(n904), .B(n885), .C(n916), .D(n894), .E(n2269), 
        .Z(n2267) );
  HS65_LL_NOR4ABX2 U10649 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .Z(
        n1136) );
  HS65_LL_AO212X4 U10650 ( .A(n863), .B(n844), .C(n875), .D(n853), .E(n1141), 
        .Z(n1139) );
  HS65_LL_NOR4ABX2 U10651 ( .A(n1513), .B(n1514), .C(n1515), .D(n1516), .Z(
        n1512) );
  HS65_LL_AO212X4 U10652 ( .A(n822), .B(n803), .C(n834), .D(n812), .E(n1517), 
        .Z(n1515) );
  HS65_LL_NOR4ABX2 U10653 ( .A(n1889), .B(n1890), .C(n1891), .D(n1892), .Z(
        n1888) );
  HS65_LL_AO212X4 U10654 ( .A(n781), .B(n762), .C(n793), .D(n771), .E(n1893), 
        .Z(n1891) );
  HS65_LL_NOR2X6 U10655 ( .A(n853), .B(n844), .Z(n1368) );
  HS65_LL_NOR3AX2 U10656 ( .A(n4908), .B(n4581), .C(n4909), .Z(n4902) );
  HS65_LL_NOR3AX2 U10657 ( .A(n4961), .B(n4598), .C(n4962), .Z(n4955) );
  HS65_LL_NOR3AX2 U10658 ( .A(n6554), .B(n6191), .C(n6555), .Z(n6548) );
  HS65_LL_NOR3AX2 U10659 ( .A(n6501), .B(n6174), .C(n6502), .Z(n6495) );
  HS65_LL_NOR3AX2 U10660 ( .A(n6403), .B(n6427), .C(n6212), .Z(n6721) );
  HS65_LL_NOR3AX2 U10661 ( .A(n4810), .B(n4834), .C(n4619), .Z(n5129) );
  HS65_LL_NOR3AX2 U10662 ( .A(n6478), .B(n6502), .C(n6320), .Z(n6839) );
  HS65_LL_NOR3AX2 U10663 ( .A(n4885), .B(n4909), .C(n4740), .Z(n5247) );
  HS65_LL_NOR3AX2 U10664 ( .A(n4938), .B(n4962), .C(n4766), .Z(n5362) );
  HS65_LL_NOR3AX2 U10665 ( .A(n6531), .B(n6555), .C(n6359), .Z(n6954) );
  HS65_LL_NOR3AX2 U10666 ( .A(n6532), .B(n6361), .C(n6192), .Z(n6528) );
  HS65_LL_NOR3AX2 U10667 ( .A(n4939), .B(n4768), .C(n4599), .Z(n4935) );
  HS65_LL_NOR3AX2 U10668 ( .A(n4695), .B(n4472), .C(n4696), .Z(n4689) );
  HS65_LL_NOR3AX2 U10669 ( .A(n6288), .B(n6065), .C(n6289), .Z(n6282) );
  HS65_LL_NAND2X7 U10670 ( .A(n419), .B(n435), .Z(n3868) );
  HS65_LL_NAND2X7 U10671 ( .A(n191), .B(n223), .Z(n3514) );
  HS65_LL_NAND2X7 U10672 ( .A(n637), .B(n648), .Z(n3753) );
  HS65_LL_NAND2X7 U10673 ( .A(n326), .B(n348), .Z(n8053) );
  HS65_LL_NOR4ABX2 U10674 ( .A(n6675), .B(n6655), .C(n6663), .D(n6632), .Z(
        n7254) );
  HS65_LL_NOR4ABX2 U10675 ( .A(n5082), .B(n5062), .C(n5070), .D(n5039), .Z(
        n5662) );
  HS65_LL_NAND2X7 U10676 ( .A(n105), .B(n125), .Z(n8830) );
  HS65_LL_NAND2X7 U10677 ( .A(n585), .B(n605), .Z(n8740) );
  HS65_LL_NAND2X7 U10678 ( .A(n110), .B(n123), .Z(n8766) );
  HS65_LL_NAND2X7 U10679 ( .A(n349), .B(n319), .Z(n8054) );
  HS65_LL_NAND2X7 U10680 ( .A(n372), .B(n387), .Z(n7985) );
  HS65_LL_NOR3AX2 U10681 ( .A(n1699), .B(n1564), .C(n1734), .Z(n1825) );
  HS65_LL_NOR3AX2 U10682 ( .A(n1323), .B(n1188), .C(n1358), .Z(n1449) );
  HS65_LL_NOR3AX2 U10683 ( .A(n2075), .B(n1940), .C(n2110), .Z(n2201) );
  HS65_LL_NOR4ABX2 U10684 ( .A(n3837), .B(n3838), .C(n3839), .D(n3840), .Z(
        n3836) );
  HS65_LL_NOR4ABX2 U10685 ( .A(n5335), .B(n5336), .C(n5337), .D(n5338), .Z(
        n4908) );
  HS65_LL_NAND3AX6 U10686 ( .A(n5339), .B(n5340), .C(n5341), .Z(n5337) );
  HS65_LL_MX41X7 U10687 ( .D0(n244), .S0(n267), .D1(n253), .S1(n236), .D2(n258), .S2(n243), .D3(n263), .S3(n237), .Z(n5338) );
  HS65_LL_NOR4ABX2 U10688 ( .A(n5347), .B(n5348), .C(n5349), .D(n5350), .Z(
        n5335) );
  HS65_LL_NOR4ABX2 U10689 ( .A(n5450), .B(n5451), .C(n5452), .D(n5453), .Z(
        n4961) );
  HS65_LL_NAND3AX6 U10690 ( .A(n5454), .B(n5455), .C(n5456), .Z(n5452) );
  HS65_LL_MX41X7 U10691 ( .D0(n461), .S0(n484), .D1(n470), .S1(n453), .D2(n475), .S2(n460), .D3(n480), .S3(n454), .Z(n5453) );
  HS65_LL_NOR4ABX2 U10692 ( .A(n5462), .B(n5463), .C(n5464), .D(n5465), .Z(
        n5450) );
  HS65_LL_NOR4ABX2 U10693 ( .A(n7042), .B(n7043), .C(n7044), .D(n7045), .Z(
        n6554) );
  HS65_LL_NAND3AX6 U10694 ( .A(n7046), .B(n7047), .C(n7048), .Z(n7044) );
  HS65_LL_MX41X7 U10695 ( .D0(n286), .S0(n309), .D1(n295), .S1(n278), .D2(n300), .S2(n285), .D3(n305), .S3(n279), .Z(n7045) );
  HS65_LL_NOR4ABX2 U10696 ( .A(n7054), .B(n7055), .C(n7056), .D(n7057), .Z(
        n7042) );
  HS65_LL_NOR4ABX2 U10697 ( .A(n6927), .B(n6928), .C(n6929), .D(n6930), .Z(
        n6501) );
  HS65_LL_NAND3AX6 U10698 ( .A(n6931), .B(n6932), .C(n6933), .Z(n6929) );
  HS65_LL_MX41X7 U10699 ( .D0(n55), .S0(n81), .D1(n88), .S1(n59), .D2(n73), 
        .S2(n56), .D3(n86), .S3(n58), .Z(n6930) );
  HS65_LL_NOR4ABX2 U10700 ( .A(n6939), .B(n6940), .C(n6941), .D(n6942), .Z(
        n6927) );
  HS65_LL_NOR4ABX2 U10701 ( .A(n1685), .B(n1686), .C(n1687), .D(n1688), .Z(
        n1684) );
  HS65_LL_NOR4ABX2 U10702 ( .A(n2483), .B(n2426), .C(n2359), .D(n2464), .Z(
        n2570) );
  HS65_LL_NOR3AX2 U10703 ( .A(n2451), .B(n2316), .C(n2486), .Z(n2577) );
  HS65_LL_NOR4ABX2 U10704 ( .A(n2100), .B(n2055), .C(n2072), .D(n2091), .Z(
        n2189) );
  HS65_LL_NAND4ABX3 U10705 ( .A(n9022), .B(n9023), .C(n9024), .D(n9025), .Z(
        n7697) );
  HS65_LL_AOI222X2 U10706 ( .A(n584), .B(n615), .C(n586), .D(n605), .E(n590), 
        .F(n616), .Z(n9024) );
  HS65_LL_NAND4ABX3 U10707 ( .A(n8151), .B(n8728), .C(n8683), .D(n8392), .Z(
        n9023) );
  HS65_LL_NOR4ABX2 U10708 ( .A(n8718), .B(n8711), .C(n8750), .D(n8695), .Z(
        n9025) );
  HS65_LL_NAND4ABX3 U10709 ( .A(n9080), .B(n9081), .C(n9082), .D(n9083), .Z(
        n7735) );
  HS65_LL_AOI222X2 U10710 ( .A(n104), .B(n135), .C(n106), .D(n125), .E(n110), 
        .F(n136), .Z(n9082) );
  HS65_LL_NAND4ABX3 U10711 ( .A(n8174), .B(n8818), .C(n8773), .D(n8444), .Z(
        n9081) );
  HS65_LL_NOR4ABX2 U10712 ( .A(n8808), .B(n8801), .C(n8840), .D(n8785), .Z(
        n9083) );
  HS65_LL_NOR4ABX2 U10713 ( .A(n3882), .B(n3827), .C(n3378), .D(n3863), .Z(
        n4305) );
  HS65_LL_NOR4ABX2 U10714 ( .A(n1348), .B(n1303), .C(n1320), .D(n1339), .Z(
        n1437) );
  HS65_LL_NOR4ABX2 U10715 ( .A(n1724), .B(n1679), .C(n1696), .D(n1715), .Z(
        n1813) );
  HS65_LL_NOR4ABX2 U10716 ( .A(n5550), .B(n5551), .C(n5552), .D(n5553), .Z(
        n5549) );
  HS65_LL_MX41X7 U10717 ( .D0(n458), .S0(n482), .D1(n457), .S1(n479), .D2(n475), .S2(n451), .D3(n450), .S3(n467), .Z(n5552) );
  HS65_LL_NOR4ABX2 U10718 ( .A(n5528), .B(n5529), .C(n5530), .D(n5531), .Z(
        n5527) );
  HS65_LL_MX41X7 U10719 ( .D0(n241), .S0(n265), .D1(n240), .S1(n262), .D2(n258), .S2(n234), .D3(n233), .S3(n250), .Z(n5530) );
  HS65_LL_NOR4ABX2 U10720 ( .A(n7142), .B(n7143), .C(n7144), .D(n7145), .Z(
        n7141) );
  HS65_LL_MX41X7 U10721 ( .D0(n283), .S0(n307), .D1(n282), .S1(n304), .D2(n300), .S2(n276), .D3(n275), .S3(n292), .Z(n7144) );
  HS65_LL_NOR4ABX2 U10722 ( .A(n7654), .B(n7717), .C(n9062), .D(n7736), .Z(
        n9061) );
  HS65_LL_MX41X7 U10723 ( .D0(n131), .S0(n99), .D1(n126), .S1(n110), .D2(n135), 
        .S2(n105), .D3(n106), .S3(n123), .Z(n9062) );
  HS65_LL_NOR4ABX2 U10724 ( .A(n5674), .B(n5568), .C(n5783), .D(n5694), .Z(
        n5782) );
  HS65_LL_MX41X7 U10725 ( .D0(n669), .S0(n695), .D1(n676), .S1(n691), .D2(n684), .S2(n679), .D3(n678), .S3(n701), .Z(n5783) );
  HS65_LL_NOR4ABX2 U10726 ( .A(n7634), .B(n7679), .C(n9004), .D(n7698), .Z(
        n9003) );
  HS65_LL_MX41X7 U10727 ( .D0(n611), .S0(n579), .D1(n606), .S1(n590), .D2(n615), .S2(n585), .D3(n586), .S3(n603), .Z(n9004) );
  HS65_LL_NOR4ABX2 U10728 ( .A(n7266), .B(n7160), .C(n7375), .D(n7286), .Z(
        n7374) );
  HS65_LL_MX41X7 U10729 ( .D0(n493), .S0(n519), .D1(n500), .S1(n515), .D2(n508), .S2(n503), .D3(n502), .S3(n525), .Z(n7375) );
  HS65_LL_NOR4ABX2 U10730 ( .A(n7120), .B(n7121), .C(n7122), .D(n7123), .Z(
        n7119) );
  HS65_LL_MX41X7 U10731 ( .D0(n57), .S0(n79), .D1(n62), .S1(n84), .D2(n73), 
        .S2(n63), .D3(n64), .S3(n91), .Z(n7122) );
  HS65_LL_NOR4ABX2 U10732 ( .A(n5644), .B(n5504), .C(n5721), .D(n5664), .Z(
        n5720) );
  HS65_LL_MX41X7 U10733 ( .D0(n14), .S0(n40), .D1(n21), .S1(n36), .D2(n24), 
        .S2(n29), .D3(n23), .S3(n46), .Z(n5721) );
  HS65_LL_NOR4ABX2 U10734 ( .A(n7236), .B(n7096), .C(n7313), .D(n7256), .Z(
        n7312) );
  HS65_LL_MX41X7 U10735 ( .D0(n536), .S0(n562), .D1(n543), .S1(n558), .D2(n546), .S2(n551), .D3(n545), .S3(n568), .Z(n7313) );
  HS65_LL_NAND2X7 U10736 ( .A(n389), .B(n372), .Z(n8271) );
  HS65_LL_NOR4ABX2 U10737 ( .A(n3447), .B(n2950), .C(n3089), .D(n3470), .Z(
        n4194) );
  HS65_LL_NAND2X7 U10738 ( .A(n132), .B(n113), .Z(n8841) );
  HS65_LL_NAND3X5 U10739 ( .A(n8946), .B(n8947), .C(n8948), .Z(n8644) );
  HS65_LL_NOR4ABX2 U10740 ( .A(n8099), .B(n8211), .C(n8112), .D(n8075), .Z(
        n8947) );
  HS65_LL_NOR4ABX2 U10741 ( .A(n8235), .B(n7853), .C(n8247), .D(n8297), .Z(
        n8946) );
  HS65_LL_NOR4ABX2 U10742 ( .A(n8285), .B(n7985), .C(n8949), .D(n8950), .Z(
        n8948) );
  HS65_LL_NOR4ABX2 U10743 ( .A(n6914), .B(n6915), .C(n6916), .D(n6917), .Z(
        n6479) );
  HS65_LL_NAND3AX6 U10744 ( .A(n6918), .B(n6919), .C(n6920), .Z(n6917) );
  HS65_LL_NAND4ABX3 U10745 ( .A(n6921), .B(n6922), .C(n6923), .D(n6924), .Z(
        n6916) );
  HS65_LL_AOI222X2 U10746 ( .A(n69), .B(n82), .C(n76), .D(n6346), .E(n68), .F(
        n77), .Z(n6914) );
  HS65_LL_NOR4ABX2 U10747 ( .A(n5280), .B(n5281), .C(n5282), .D(n5283), .Z(
        n5274) );
  HS65_LL_NOR4ABX2 U10748 ( .A(n6872), .B(n6873), .C(n6874), .D(n6875), .Z(
        n6866) );
  HS65_LL_NOR4ABX2 U10749 ( .A(n6987), .B(n6988), .C(n6989), .D(n6990), .Z(
        n6981) );
  HS65_LL_NAND2X7 U10750 ( .A(n454), .B(n477), .Z(n5386) );
  HS65_LL_NAND2X7 U10751 ( .A(n237), .B(n260), .Z(n5271) );
  HS65_LL_NAND2X7 U10752 ( .A(n279), .B(n302), .Z(n6978) );
  HS65_LL_NAND2X7 U10753 ( .A(n58), .B(n83), .Z(n6863) );
  HS65_LL_NOR4ABX2 U10754 ( .A(n5084), .B(n5085), .C(n5086), .D(n5087), .Z(
        n4695) );
  HS65_LL_MX41X7 U10755 ( .D0(n41), .S0(n15), .D1(n45), .S1(n19), .D2(n17), 
        .S2(n29), .D3(n18), .S3(n34), .Z(n5087) );
  HS65_LL_NAND3AX6 U10756 ( .A(n5088), .B(n5089), .C(n5090), .Z(n5086) );
  HS65_LL_NOR4ABX2 U10757 ( .A(n5092), .B(n5093), .C(n5094), .D(n5095), .Z(
        n5085) );
  HS65_LL_NOR4ABX2 U10758 ( .A(n6677), .B(n6678), .C(n6679), .D(n6680), .Z(
        n6288) );
  HS65_LL_MX41X7 U10759 ( .D0(n563), .S0(n537), .D1(n567), .S1(n541), .D2(n539), .S2(n551), .D3(n540), .S3(n556), .Z(n6680) );
  HS65_LL_NAND3AX6 U10760 ( .A(n6681), .B(n6682), .C(n6683), .Z(n6679) );
  HS65_LL_NOR4ABX2 U10761 ( .A(n6685), .B(n6686), .C(n6687), .D(n6688), .Z(
        n6678) );
  HS65_LL_NOR4ABX2 U10762 ( .A(n8732), .B(n8733), .C(n8734), .D(n8735), .Z(
        n8376) );
  HS65_LL_NAND3AX6 U10763 ( .A(n8736), .B(n7808), .C(n8737), .Z(n8735) );
  HS65_LL_NAND4ABX3 U10764 ( .A(n8738), .B(n8739), .C(n8740), .D(n7794), .Z(
        n8734) );
  HS65_LL_AOI222X2 U10765 ( .A(n584), .B(n609), .C(n614), .D(n8130), .E(n583), 
        .F(n616), .Z(n8732) );
  HS65_LL_NOR4ABX2 U10766 ( .A(n3760), .B(n3716), .C(n3732), .D(n3751), .Z(
        n4241) );
  HS65_LL_NOR4ABX2 U10767 ( .A(n3322), .B(n3323), .C(n3324), .D(n3325), .Z(
        n3316) );
  HS65_LL_NAND2X7 U10768 ( .A(n353), .B(n317), .Z(n8559) );
  HS65_LL_NAND2X7 U10769 ( .A(n325), .B(n354), .Z(n8367) );
  HS65_LL_NAND2X7 U10770 ( .A(n343), .B(n317), .Z(n8513) );
  HS65_LL_NOR4ABX2 U10771 ( .A(n4918), .B(n4919), .C(n4920), .D(n4921), .Z(
        n4912) );
  HS65_LL_NOR4ABX2 U10772 ( .A(n6564), .B(n6565), .C(n6566), .D(n6567), .Z(
        n6558) );
  HS65_LL_NOR4ABX2 U10773 ( .A(n6511), .B(n6512), .C(n6513), .D(n6514), .Z(
        n6505) );
  HS65_LL_NAND2X7 U10774 ( .A(n460), .B(n469), .Z(n5358) );
  HS65_LL_NAND2X7 U10775 ( .A(n285), .B(n294), .Z(n6950) );
  HS65_LL_NAND2X7 U10776 ( .A(n243), .B(n252), .Z(n5243) );
  HS65_LL_NAND2X7 U10777 ( .A(n56), .B(n89), .Z(n6835) );
  HS65_LL_NAND2X7 U10778 ( .A(n672), .B(n702), .Z(n5125) );
  HS65_LL_NAND2X7 U10779 ( .A(n496), .B(n526), .Z(n6717) );
  HS65_LL_NAND2X7 U10780 ( .A(n370), .B(n383), .Z(n8197) );
  HS65_LL_NAND4ABX3 U10781 ( .A(n8241), .B(n8242), .C(n8243), .D(n8244), .Z(
        n7973) );
  HS65_LL_NAND4ABX3 U10782 ( .A(n8255), .B(n8256), .C(n8257), .D(n7744), .Z(
        n8241) );
  HS65_LL_NOR3AX2 U10783 ( .A(n8249), .B(n8250), .C(n8251), .Z(n8243) );
  HS65_LL_NOR4ABX2 U10784 ( .A(n8245), .B(n8246), .C(n8247), .D(n8248), .Z(
        n8244) );
  HS65_LL_NAND2X7 U10785 ( .A(n580), .B(n602), .Z(n8669) );
  HS65_LL_NAND2X7 U10786 ( .A(n100), .B(n122), .Z(n8759) );
  HS65_LL_NAND4ABX3 U10787 ( .A(n3718), .B(n3719), .C(n3720), .D(n3721), .Z(
        n3143) );
  HS65_LL_NAND4ABX3 U10788 ( .A(n3732), .B(n3733), .C(n3734), .D(n3735), .Z(
        n3718) );
  HS65_LL_NOR3AX2 U10789 ( .A(n3726), .B(n3727), .C(n3728), .Z(n3720) );
  HS65_LL_NOR4ABX2 U10790 ( .A(n3722), .B(n3723), .C(n3724), .D(n3725), .Z(
        n3721) );
  HS65_LL_NAND4ABX3 U10791 ( .A(n8678), .B(n8679), .C(n8680), .D(n8681), .Z(
        n8138) );
  HS65_LL_NOR4ABX2 U10792 ( .A(n8682), .B(n8683), .C(n7691), .D(n7789), .Z(
        n8681) );
  HS65_LL_NOR3AX2 U10793 ( .A(n8684), .B(n7829), .C(n8685), .Z(n8680) );
  HS65_LL_NAND4ABX3 U10794 ( .A(n7672), .B(n8689), .C(n8690), .D(n7809), .Z(
        n8678) );
  HS65_LL_NAND4ABX3 U10795 ( .A(n8768), .B(n8769), .C(n8770), .D(n8771), .Z(
        n8161) );
  HS65_LL_NOR4ABX2 U10796 ( .A(n8772), .B(n8773), .C(n7729), .D(n7888), .Z(
        n8771) );
  HS65_LL_NOR3AX2 U10797 ( .A(n8774), .B(n7927), .C(n8775), .Z(n8770) );
  HS65_LL_NAND4ABX3 U10798 ( .A(n7710), .B(n8779), .C(n8780), .D(n7907), .Z(
        n8768) );
  HS65_LL_IVX9 U10799 ( .A(n2830), .Z(n411) );
  HS65_LL_NAND2X7 U10800 ( .A(n54), .B(n89), .Z(n6862) );
  HS65_LL_NAND2X7 U10801 ( .A(n96), .B(n122), .Z(n8780) );
  HS65_LL_NAND2X7 U10802 ( .A(n576), .B(n602), .Z(n8690) );
  HS65_LL_NAND2X7 U10803 ( .A(n823), .B(n812), .Z(n1718) );
  HS65_LL_NAND2X7 U10804 ( .A(n864), .B(n853), .Z(n1342) );
  HS65_LL_NAND2X7 U10805 ( .A(n782), .B(n771), .Z(n2094) );
  HS65_LL_NAND2X7 U10806 ( .A(n245), .B(n257), .Z(n5289) );
  HS65_LL_NAND2X7 U10807 ( .A(n69), .B(n76), .Z(n6881) );
  HS65_LL_NAND2X7 U10808 ( .A(n905), .B(n894), .Z(n2470) );
  HS65_LL_NAND2X7 U10809 ( .A(n419), .B(n432), .Z(n3869) );
  HS65_LL_NAND2X7 U10810 ( .A(n637), .B(n645), .Z(n3754) );
  HS65_LL_NAND4ABX3 U10811 ( .A(n2186), .B(n2187), .C(n2188), .D(n2189), .Z(
        n2131) );
  HS65_LL_NAND4ABX3 U10812 ( .A(n2002), .B(n1968), .C(n1942), .D(n1981), .Z(
        n2187) );
  HS65_LL_NAND4ABX3 U10813 ( .A(n2123), .B(n2039), .C(n2026), .D(n2190), .Z(
        n2186) );
  HS65_LL_AOI222X2 U10814 ( .A(n758), .B(n786), .C(n770), .D(n790), .E(n772), 
        .F(n785), .Z(n2188) );
  HS65_LL_NAND4ABX3 U10815 ( .A(n1815), .B(n1816), .C(n1817), .D(n1818), .Z(
        n1500) );
  HS65_LL_AOI222X2 U10816 ( .A(n821), .B(n798), .C(n801), .D(n825), .E(n834), 
        .F(n812), .Z(n1817) );
  HS65_LL_NOR4ABX2 U10817 ( .A(n1731), .B(n1674), .C(n1607), .D(n1712), .Z(
        n1818) );
  HS65_LL_NAND4ABX3 U10818 ( .A(n1689), .B(n1567), .C(n1617), .D(n1666), .Z(
        n1816) );
  HS65_LL_NAND4ABX3 U10819 ( .A(n1434), .B(n1435), .C(n1436), .D(n1437), .Z(
        n1379) );
  HS65_LL_NAND4ABX3 U10820 ( .A(n1250), .B(n1216), .C(n1190), .D(n1229), .Z(
        n1435) );
  HS65_LL_NAND4ABX3 U10821 ( .A(n1371), .B(n1287), .C(n1274), .D(n1438), .Z(
        n1434) );
  HS65_LL_AOI222X2 U10822 ( .A(n840), .B(n868), .C(n852), .D(n872), .E(n854), 
        .F(n867), .Z(n1436) );
  HS65_LL_NAND4ABX3 U10823 ( .A(n1810), .B(n1811), .C(n1812), .D(n1813), .Z(
        n1755) );
  HS65_LL_NAND4ABX3 U10824 ( .A(n1626), .B(n1592), .C(n1566), .D(n1605), .Z(
        n1811) );
  HS65_LL_NAND4ABX3 U10825 ( .A(n1747), .B(n1663), .C(n1650), .D(n1814), .Z(
        n1810) );
  HS65_LL_AOI222X2 U10826 ( .A(n799), .B(n827), .C(n811), .D(n831), .E(n813), 
        .F(n826), .Z(n1812) );
  HS65_LL_NAND4ABX3 U10827 ( .A(n2562), .B(n2563), .C(n2564), .D(n2565), .Z(
        n2507) );
  HS65_LL_NAND4ABX3 U10828 ( .A(n2378), .B(n2344), .C(n2318), .D(n2357), .Z(
        n2563) );
  HS65_LL_NAND4ABX3 U10829 ( .A(n2499), .B(n2415), .C(n2402), .D(n2566), .Z(
        n2562) );
  HS65_LL_NOR4ABX2 U10830 ( .A(n2476), .B(n2431), .C(n2448), .D(n2467), .Z(
        n2565) );
  HS65_LL_NAND4ABX3 U10831 ( .A(n1439), .B(n1440), .C(n1441), .D(n1442), .Z(
        n1124) );
  HS65_LL_AOI222X2 U10832 ( .A(n862), .B(n839), .C(n842), .D(n866), .E(n875), 
        .F(n853), .Z(n1441) );
  HS65_LL_NOR4ABX2 U10833 ( .A(n1355), .B(n1298), .C(n1231), .D(n1336), .Z(
        n1442) );
  HS65_LL_NAND4ABX3 U10834 ( .A(n1313), .B(n1191), .C(n1241), .D(n1290), .Z(
        n1440) );
  HS65_LL_NAND4ABX3 U10835 ( .A(n2191), .B(n2192), .C(n2193), .D(n2194), .Z(
        n1876) );
  HS65_LL_AOI222X2 U10836 ( .A(n780), .B(n757), .C(n760), .D(n784), .E(n793), 
        .F(n771), .Z(n2193) );
  HS65_LL_NAND4ABX3 U10837 ( .A(n2065), .B(n1943), .C(n1993), .D(n2042), .Z(
        n2192) );
  HS65_LL_NOR4ABX2 U10838 ( .A(n2107), .B(n2050), .C(n1983), .D(n2088), .Z(
        n2194) );
  HS65_LL_NAND4ABX3 U10839 ( .A(n2567), .B(n2568), .C(n2569), .D(n2570), .Z(
        n2252) );
  HS65_LL_AOI222X2 U10840 ( .A(n903), .B(n880), .C(n883), .D(n907), .E(n916), 
        .F(n894), .Z(n2569) );
  HS65_LL_NAND4ABX3 U10841 ( .A(n2441), .B(n2319), .C(n2369), .D(n2418), .Z(
        n2568) );
  HS65_LL_NAND4ABX3 U10842 ( .A(n2404), .B(n2500), .C(n2571), .D(n2379), .Z(
        n2567) );
  HS65_LL_IVX9 U10843 ( .A(n7952), .Z(n327) );
  HS65_LL_NAND2X7 U10844 ( .A(n351), .B(n334), .Z(n8347) );
  HS65_LL_NAND2X7 U10845 ( .A(n317), .B(n345), .Z(n8341) );
  HS65_LL_NAND2X7 U10846 ( .A(n377), .B(n393), .Z(n7744) );
  HS65_LL_NAND2X7 U10847 ( .A(n637), .B(n646), .Z(n3322) );
  HS65_LL_NAND2X7 U10848 ( .A(n913), .B(n885), .Z(n2397) );
  HS65_LL_NAND2X7 U10849 ( .A(n790), .B(n762), .Z(n2021) );
  HS65_LL_NAND2X7 U10850 ( .A(n872), .B(n844), .Z(n1269) );
  HS65_LL_NAND2X7 U10851 ( .A(n23), .B(n33), .Z(n5092) );
  HS65_LL_NAND2X7 U10852 ( .A(n545), .B(n555), .Z(n6685) );
  HS65_LL_NAND2X7 U10853 ( .A(n831), .B(n803), .Z(n1645) );
  HS65_LL_IVX9 U10854 ( .A(n7869), .Z(n106) );
  HS65_LL_IVX9 U10855 ( .A(n7806), .Z(n586) );
  HS65_LL_NAND2X7 U10856 ( .A(n629), .B(n650), .Z(n3669) );
  HS65_LL_NAND2X7 U10857 ( .A(n630), .B(n646), .Z(n3335) );
  HS65_LL_NAND2X7 U10858 ( .A(n155), .B(n169), .Z(n3619) );
  HS65_LL_NAND2X7 U10859 ( .A(n450), .B(n474), .Z(n5458) );
  HS65_LL_NAND2X7 U10860 ( .A(n275), .B(n299), .Z(n7050) );
  HS65_LL_NAND2X7 U10861 ( .A(n233), .B(n257), .Z(n5343) );
  HS65_LL_NAND2X7 U10862 ( .A(n64), .B(n76), .Z(n6935) );
  HS65_LL_NAND2X7 U10863 ( .A(n678), .B(n688), .Z(n5228) );
  HS65_LL_NAND2X7 U10864 ( .A(n502), .B(n512), .Z(n6820) );
  HS65_LL_NAND2X7 U10865 ( .A(n766), .B(n785), .Z(n1919) );
  HS65_LL_NAND2X7 U10866 ( .A(n807), .B(n826), .Z(n1543) );
  HS65_LL_NAND2X7 U10867 ( .A(n848), .B(n867), .Z(n1167) );
  HS65_LL_NAND2X7 U10868 ( .A(n889), .B(n908), .Z(n2295) );
  HS65_LL_NAND2X7 U10869 ( .A(n626), .B(n646), .Z(n3716) );
  HS65_LL_NAND2X7 U10870 ( .A(n376), .B(n398), .Z(n8078) );
  HS65_LL_NAND2X7 U10871 ( .A(n411), .B(n441), .Z(n3784) );
  HS65_LL_NAND2X7 U10872 ( .A(n580), .B(n610), .Z(n8697) );
  HS65_LL_NAND2X7 U10873 ( .A(n100), .B(n130), .Z(n8787) );
  HS65_LL_IVX9 U10874 ( .A(n3005), .Z(n316) );
  HS65_LL_NAND2X7 U10875 ( .A(n149), .B(n169), .Z(n3262) );
  HS65_LL_NAND2X7 U10876 ( .A(n197), .B(n221), .Z(n3426) );
  HS65_LL_NAND2X7 U10877 ( .A(n375), .B(n393), .Z(n8220) );
  HS65_LL_NAND2X7 U10878 ( .A(n539), .B(n563), .Z(n6635) );
  HS65_LL_NAND2X7 U10879 ( .A(n17), .B(n41), .Z(n5042) );
  HS65_LL_NAND2X7 U10880 ( .A(n661), .B(n625), .Z(n3701) );
  HS65_LL_NAND2X7 U10881 ( .A(n371), .B(n390), .Z(n8286) );
  HS65_LL_NOR3X4 U10882 ( .A(n7899), .B(n7648), .C(n7718), .Z(n7865) );
  HS65_LL_NAND2X7 U10883 ( .A(n341), .B(n325), .Z(n8335) );
  HS65_LL_NAND2X7 U10884 ( .A(n576), .B(n607), .Z(n7797) );
  HS65_LL_NAND2X7 U10885 ( .A(n96), .B(n127), .Z(n7896) );
  HS65_LL_NAND2X7 U10886 ( .A(n844), .B(n867), .Z(n1348) );
  HS65_LL_NAND2X7 U10887 ( .A(n885), .B(n908), .Z(n2476) );
  HS65_LL_NAND2X7 U10888 ( .A(n762), .B(n785), .Z(n2100) );
  HS65_LL_NAND2X7 U10889 ( .A(n803), .B(n826), .Z(n1724) );
  HS65_LL_NAND2X7 U10890 ( .A(n391), .B(n374), .Z(n8102) );
  HS65_LL_NOR3X4 U10891 ( .A(n4511), .B(n4512), .C(n4513), .Z(n4488) );
  HS65_LL_NOR3X4 U10892 ( .A(n6104), .B(n6105), .C(n6106), .Z(n6081) );
  HS65_LL_NOR3X4 U10893 ( .A(n7773), .B(n8622), .C(n8623), .Z(n8611) );
  HS65_LL_NAND2X7 U10894 ( .A(n653), .B(n627), .Z(n3139) );
  HS65_LL_NAND2X7 U10895 ( .A(n240), .B(n260), .Z(n4737) );
  HS65_LL_NAND2X7 U10896 ( .A(n457), .B(n477), .Z(n4798) );
  HS65_LL_NAND2X7 U10897 ( .A(n282), .B(n302), .Z(n6391) );
  HS65_LL_NAND2X7 U10898 ( .A(n62), .B(n83), .Z(n6352) );
  HS65_LL_NAND2X7 U10899 ( .A(n500), .B(n514), .Z(n6245) );
  HS65_LL_NAND2X7 U10900 ( .A(n676), .B(n690), .Z(n4652) );
  HS65_LL_NAND3X5 U10901 ( .A(n8699), .B(n8700), .C(n8701), .Z(n8692) );
  HS65_LL_AOI12X2 U10902 ( .A(n585), .B(n599), .C(n7837), .Z(n8701) );
  HS65_LL_NAND3X5 U10903 ( .A(n8789), .B(n8790), .C(n8791), .Z(n8782) );
  HS65_LL_AOI12X2 U10904 ( .A(n105), .B(n119), .C(n7876), .Z(n8791) );
  HS65_LL_NAND2X7 U10905 ( .A(n848), .B(n871), .Z(n1310) );
  HS65_LL_NAND2X7 U10906 ( .A(n766), .B(n789), .Z(n2062) );
  HS65_LL_NAND2X7 U10907 ( .A(n436), .B(n407), .Z(n3838) );
  HS65_LL_NAND2X7 U10908 ( .A(n658), .B(n626), .Z(n3763) );
  HS65_LL_NAND2X7 U10909 ( .A(n769), .B(n785), .Z(n2099) );
  HS65_LL_NAND2X7 U10910 ( .A(n810), .B(n826), .Z(n1723) );
  HS65_LL_NAND2X7 U10911 ( .A(n892), .B(n908), .Z(n2475) );
  HS65_LL_NAND2X7 U10912 ( .A(n851), .B(n867), .Z(n1347) );
  HS65_LL_NAND2X7 U10913 ( .A(n889), .B(n912), .Z(n2438) );
  HS65_LL_NAND2X7 U10914 ( .A(n807), .B(n830), .Z(n1686) );
  HS65_LL_NAND2X7 U10915 ( .A(n88), .B(n58), .Z(n6902) );
  HS65_LL_NAND2X7 U10916 ( .A(n253), .B(n237), .Z(n5310) );
  HS65_LL_NAND2X7 U10917 ( .A(n470), .B(n454), .Z(n5425) );
  HS65_LL_NAND2X7 U10918 ( .A(n295), .B(n279), .Z(n7017) );
  HS65_LL_NAND2X7 U10919 ( .A(n389), .B(n374), .Z(n8281) );
  HS65_LL_AOI12X2 U10920 ( .A(n901), .B(n895), .C(n2478), .Z(n2477) );
  HS65_LL_AOI12X2 U10921 ( .A(n819), .B(n813), .C(n1726), .Z(n1725) );
  HS65_LL_AOI12X2 U10922 ( .A(n860), .B(n854), .C(n1350), .Z(n1349) );
  HS65_LL_AOI12X2 U10923 ( .A(n778), .B(n772), .C(n2102), .Z(n2101) );
  HS65_LL_NAND2X7 U10924 ( .A(n216), .B(n200), .Z(n3483) );
  HS65_LL_NAND2X7 U10925 ( .A(n585), .B(n607), .Z(n8708) );
  HS65_LL_NAND2X7 U10926 ( .A(n105), .B(n127), .Z(n8798) );
  HS65_LL_NAND2X7 U10927 ( .A(n580), .B(n607), .Z(n8402) );
  HS65_LL_NAND2X7 U10928 ( .A(n100), .B(n127), .Z(n8454) );
  HS65_LL_NAND2X7 U10929 ( .A(n807), .B(n832), .Z(n1618) );
  HS65_LL_NAND2X7 U10930 ( .A(n436), .B(n417), .Z(n3389) );
  HS65_LL_NAND2X7 U10931 ( .A(n216), .B(n194), .Z(n3106) );
  HS65_LL_NAND2X7 U10932 ( .A(n906), .B(n890), .Z(n2450) );
  HS65_LL_NAND2X7 U10933 ( .A(n889), .B(n914), .Z(n2370) );
  HS65_LL_AOI12X2 U10934 ( .A(n624), .B(n651), .C(n3762), .Z(n3761) );
  HS65_LL_AOI12X2 U10935 ( .A(n405), .B(n442), .C(n3877), .Z(n3876) );
  HS65_LL_AOI12X2 U10936 ( .A(n201), .B(n219), .C(n3523), .Z(n3522) );
  HS65_LL_NAND2X7 U10937 ( .A(n766), .B(n791), .Z(n1994) );
  HS65_LL_NAND2X7 U10938 ( .A(n848), .B(n873), .Z(n1242) );
  HS65_LL_NAND3AX6 U10939 ( .A(n1610), .B(n1611), .C(n1612), .Z(n1597) );
  HS65_LL_AOI12X2 U10940 ( .A(n827), .B(n1613), .C(n1614), .Z(n1612) );
  HS65_LL_NAND2X7 U10941 ( .A(n783), .B(n767), .Z(n2074) );
  HS65_LL_NAND2X7 U10942 ( .A(n865), .B(n849), .Z(n1322) );
  HS65_LL_IVX9 U10943 ( .A(n2775), .Z(n574) );
  HS65_LL_NAND3X5 U10944 ( .A(n5915), .B(n5916), .C(n5917), .Z(n5553) );
  HS65_LL_NOR4ABX2 U10945 ( .A(n5435), .B(n4944), .C(n4982), .D(n4970), .Z(
        n5916) );
  HS65_LL_NOR4ABX2 U10946 ( .A(n5376), .B(n4605), .C(n5423), .D(n5444), .Z(
        n5915) );
  HS65_LL_NOR4X4 U10947 ( .A(n5417), .B(n4786), .C(n5918), .D(n5919), .Z(n5917) );
  HS65_LL_NAND3X5 U10948 ( .A(n7507), .B(n7508), .C(n7509), .Z(n7145) );
  HS65_LL_NOR4ABX2 U10949 ( .A(n7027), .B(n6537), .C(n6575), .D(n6563), .Z(
        n7508) );
  HS65_LL_NOR4ABX2 U10950 ( .A(n6968), .B(n6198), .C(n7015), .D(n7036), .Z(
        n7507) );
  HS65_LL_NOR4X4 U10951 ( .A(n7009), .B(n6379), .C(n7510), .D(n7511), .Z(n7509) );
  HS65_LL_NAND3X5 U10952 ( .A(n5856), .B(n5857), .C(n5858), .Z(n5531) );
  HS65_LL_NOR4ABX2 U10953 ( .A(n5320), .B(n4891), .C(n4929), .D(n4917), .Z(
        n5857) );
  HS65_LL_NOR4ABX2 U10954 ( .A(n5261), .B(n4588), .C(n5308), .D(n5329), .Z(
        n5856) );
  HS65_LL_NOR4X4 U10955 ( .A(n5302), .B(n4759), .C(n5859), .D(n5860), .Z(n5858) );
  HS65_LL_NAND3X5 U10956 ( .A(n7448), .B(n7449), .C(n7450), .Z(n7123) );
  HS65_LL_NOR4ABX2 U10957 ( .A(n6912), .B(n6484), .C(n6522), .D(n6510), .Z(
        n7449) );
  HS65_LL_NOR4ABX2 U10958 ( .A(n6853), .B(n6181), .C(n6900), .D(n6921), .Z(
        n7448) );
  HS65_LL_NOR4X4 U10959 ( .A(n6894), .B(n6340), .C(n7451), .D(n7452), .Z(n7450) );
  HS65_LL_NAND3X5 U10960 ( .A(n5784), .B(n5785), .C(n5786), .Z(n5694) );
  HS65_LL_NOR4ABX2 U10961 ( .A(n5204), .B(n4816), .C(n4856), .D(n4842), .Z(
        n5785) );
  HS65_LL_NOR4ABX2 U10962 ( .A(n5144), .B(n4536), .C(n5192), .D(n5213), .Z(
        n5784) );
  HS65_LL_NOR4X4 U10963 ( .A(n5186), .B(n4640), .C(n5787), .D(n5788), .Z(n5786) );
  HS65_LL_NAND3X5 U10964 ( .A(n7376), .B(n7377), .C(n7378), .Z(n7286) );
  HS65_LL_NOR4ABX2 U10965 ( .A(n6796), .B(n6409), .C(n6449), .D(n6435), .Z(
        n7377) );
  HS65_LL_NOR4ABX2 U10966 ( .A(n6736), .B(n6129), .C(n6784), .D(n6805), .Z(
        n7376) );
  HS65_LL_NOR4X4 U10967 ( .A(n6778), .B(n6233), .C(n7379), .D(n7380), .Z(n7378) );
  HS65_LL_NAND2X7 U10968 ( .A(n824), .B(n808), .Z(n1698) );
  HS65_LL_NAND2X7 U10969 ( .A(n107), .B(n131), .Z(n8827) );
  HS65_LL_NAND2X7 U10970 ( .A(n587), .B(n611), .Z(n8737) );
  HS65_LL_NAND2X7 U10971 ( .A(n415), .B(n440), .Z(n3849) );
  HS65_LL_AOI12X2 U10972 ( .A(n592), .B(n616), .C(n8710), .Z(n8709) );
  HS65_LL_AOI12X2 U10973 ( .A(n112), .B(n136), .C(n8800), .Z(n8799) );
  HS65_LL_NAND2X7 U10974 ( .A(n592), .B(n611), .Z(n7670) );
  HS65_LL_NAND3X5 U10975 ( .A(n7314), .B(n7315), .C(n7316), .Z(n7256) );
  HS65_LL_NOR4ABX2 U10976 ( .A(n6664), .B(n6073), .C(n6616), .D(n6700), .Z(
        n7314) );
  HS65_LL_NOR4ABX2 U10977 ( .A(n6673), .B(n6270), .C(n6311), .D(n6297), .Z(
        n7315) );
  HS65_LL_NOR4X4 U10978 ( .A(n6657), .B(n6156), .C(n7317), .D(n7318), .Z(n7316) );
  HS65_LL_NAND3X5 U10979 ( .A(n5722), .B(n5723), .C(n5724), .Z(n5664) );
  HS65_LL_NOR4ABX2 U10980 ( .A(n5071), .B(n4480), .C(n5023), .D(n5107), .Z(
        n5722) );
  HS65_LL_NOR4ABX2 U10981 ( .A(n5080), .B(n4677), .C(n4718), .D(n4704), .Z(
        n5723) );
  HS65_LL_NOR4X4 U10982 ( .A(n5064), .B(n4563), .C(n5725), .D(n5726), .Z(n5724) );
  HS65_LL_NAND2X7 U10983 ( .A(n393), .B(n374), .Z(n8282) );
  HS65_LL_NAND2X7 U10984 ( .A(n633), .B(n649), .Z(n3734) );
  HS65_LL_OAI21X3 U10985 ( .A(n460), .B(n458), .C(n472), .Z(n5932) );
  HS65_LL_OAI21X3 U10986 ( .A(n285), .B(n283), .C(n297), .Z(n7524) );
  HS65_LL_OAI21X3 U10987 ( .A(n243), .B(n241), .C(n255), .Z(n5873) );
  HS65_LL_OAI21X3 U10988 ( .A(n56), .B(n57), .C(n90), .Z(n7467) );
  HS65_LL_OAI21X3 U10989 ( .A(n496), .B(n493), .C(n523), .Z(n7358) );
  HS65_LL_NAND2X7 U10990 ( .A(n847), .B(n871), .Z(n1351) );
  HS65_LL_NAND2X7 U10991 ( .A(n765), .B(n789), .Z(n2103) );
  HS65_LL_NAND2X7 U10992 ( .A(n629), .B(n660), .Z(n3298) );
  HS65_LL_NAND2X7 U10993 ( .A(n788), .B(n763), .Z(n1935) );
  HS65_LL_NAND2X7 U10994 ( .A(n870), .B(n845), .Z(n1183) );
  HS65_LL_NAND2X7 U10995 ( .A(n427), .B(n407), .Z(n3878) );
  HS65_LL_NAND2X7 U10996 ( .A(n813), .B(n832), .Z(n1602) );
  HS65_LL_NAND2X7 U10997 ( .A(n810), .B(n832), .Z(n1714) );
  HS65_LL_NAND2X7 U10998 ( .A(n636), .B(n653), .Z(n3749) );
  HS65_LL_NAND2X7 U10999 ( .A(n428), .B(n417), .Z(n3865) );
  HS65_LL_NAND2X7 U11000 ( .A(n442), .B(n417), .Z(n3373) );
  HS65_LL_NAND2X7 U11001 ( .A(n212), .B(n194), .Z(n3511) );
  HS65_LL_NAND2X7 U11002 ( .A(n219), .B(n194), .Z(n3088) );
  HS65_LL_NAND2X7 U11003 ( .A(n911), .B(n886), .Z(n2311) );
  HS65_LL_NAND2X7 U11004 ( .A(n903), .B(n890), .Z(n2402) );
  HS65_LL_IVX9 U11005 ( .A(n2749), .Z(n404) );
  HS65_LL_NAND2X7 U11006 ( .A(n895), .B(n914), .Z(n2354) );
  HS65_LL_NAND2X7 U11007 ( .A(n892), .B(n914), .Z(n2466) );
  HS65_LL_NAND2X7 U11008 ( .A(n772), .B(n791), .Z(n1978) );
  HS65_LL_NAND2X7 U11009 ( .A(n854), .B(n873), .Z(n1226) );
  HS65_LL_NAND2X7 U11010 ( .A(n851), .B(n873), .Z(n1338) );
  HS65_LL_NAND2X7 U11011 ( .A(n769), .B(n791), .Z(n2090) );
  HS65_LL_NAND2X7 U11012 ( .A(n888), .B(n912), .Z(n2479) );
  HS65_LL_NAND2X7 U11013 ( .A(n806), .B(n830), .Z(n1727) );
  HS65_LL_NAND2X7 U11014 ( .A(n780), .B(n767), .Z(n2026) );
  HS65_LL_NAND2X7 U11015 ( .A(n862), .B(n849), .Z(n1274) );
  HS65_LL_NAND2X7 U11016 ( .A(n66), .B(n79), .Z(n6920) );
  HS65_LL_NAND2X7 U11017 ( .A(n235), .B(n265), .Z(n5328) );
  HS65_LL_NAND2X7 U11018 ( .A(n452), .B(n482), .Z(n5443) );
  HS65_LL_NAND2X7 U11019 ( .A(n680), .B(n695), .Z(n5212) );
  HS65_LL_NAND2X7 U11020 ( .A(n25), .B(n40), .Z(n5106) );
  HS65_LL_NAND2X7 U11021 ( .A(n277), .B(n307), .Z(n7035) );
  HS65_LL_NAND2X7 U11022 ( .A(n504), .B(n519), .Z(n6804) );
  HS65_LL_NAND2X7 U11023 ( .A(n547), .B(n562), .Z(n6699) );
  HS65_LL_NAND2X7 U11024 ( .A(n821), .B(n808), .Z(n1650) );
  HS65_LL_NAND2X7 U11025 ( .A(n209), .B(n200), .Z(n3524) );
  HS65_LL_NAND2X7 U11026 ( .A(n566), .B(n532), .Z(n6073) );
  HS65_LL_NAND2X7 U11027 ( .A(n44), .B(n10), .Z(n4480) );
  HS65_LL_NAND2X7 U11028 ( .A(n834), .B(n814), .Z(n1611) );
  HS65_LL_NAND2X7 U11029 ( .A(n916), .B(n896), .Z(n2363) );
  HS65_LL_NAND2X7 U11030 ( .A(n875), .B(n855), .Z(n1235) );
  HS65_LL_NAND2X7 U11031 ( .A(n651), .B(n635), .Z(n3319) );
  HS65_LL_NAND2X7 U11032 ( .A(n793), .B(n773), .Z(n1987) );
  HS65_LL_NAND2X7 U11033 ( .A(n355), .B(n325), .Z(n8584) );
  HS65_LL_NAND2X7 U11034 ( .A(n340), .B(n334), .Z(n8569) );
  HS65_LL_NAND2X7 U11035 ( .A(n639), .B(n649), .Z(n3674) );
  HS65_LL_NAND2X7 U11036 ( .A(n523), .B(n490), .Z(n6129) );
  HS65_LL_NAND2X7 U11037 ( .A(n699), .B(n666), .Z(n4536) );
  HS65_LL_NAND2X7 U11038 ( .A(n255), .B(n247), .Z(n4588) );
  HS65_LL_NAND2X7 U11039 ( .A(n297), .B(n289), .Z(n6198) );
  HS65_LL_NAND2X7 U11040 ( .A(n90), .B(n68), .Z(n6181) );
  HS65_LL_NAND2X7 U11041 ( .A(n472), .B(n464), .Z(n4605) );
  HS65_LL_NAND2X7 U11042 ( .A(n242), .B(n256), .Z(n5284) );
  HS65_LL_NAND2X7 U11043 ( .A(n54), .B(n74), .Z(n6876) );
  HS65_LL_OAI21X3 U11044 ( .A(n875), .B(n868), .C(n851), .Z(n1166) );
  HS65_LL_AOI12X2 U11045 ( .A(n261), .B(n242), .C(n5342), .Z(n5341) );
  HS65_LL_AOI12X2 U11046 ( .A(n303), .B(n284), .C(n7049), .Z(n7048) );
  HS65_LL_AOI12X2 U11047 ( .A(n85), .B(n54), .C(n6934), .Z(n6933) );
  HS65_LL_NAND2X7 U11048 ( .A(n64), .B(n79), .Z(n6474) );
  HS65_LL_NAND2X7 U11049 ( .A(n341), .B(n328), .Z(n8525) );
  HS65_LL_OAI21X3 U11050 ( .A(n539), .B(n536), .C(n566), .Z(n7296) );
  HS65_LL_OAI21X3 U11051 ( .A(n17), .B(n14), .C(n44), .Z(n5704) );
  HS65_LL_NAND2X7 U11052 ( .A(n640), .B(n660), .Z(n3328) );
  HS65_LL_NAND2X7 U11053 ( .A(n457), .B(n482), .Z(n4968) );
  HS65_LL_NAND2X7 U11054 ( .A(n282), .B(n307), .Z(n6561) );
  HS65_LL_NAND2X7 U11055 ( .A(n240), .B(n265), .Z(n4915) );
  HS65_LL_NAND2X7 U11056 ( .A(n62), .B(n79), .Z(n6508) );
  HS65_LL_NAND2X7 U11057 ( .A(n246), .B(n256), .Z(n5344) );
  HS65_LL_NAND2X7 U11058 ( .A(n463), .B(n473), .Z(n5459) );
  HS65_LL_NAND2X7 U11059 ( .A(n288), .B(n298), .Z(n7051) );
  HS65_LL_NAND2X7 U11060 ( .A(n67), .B(n74), .Z(n6936) );
  HS65_LL_NAND2X7 U11061 ( .A(n599), .B(n583), .Z(n8003) );
  HS65_LL_NAND2X7 U11062 ( .A(n119), .B(n103), .Z(n8016) );
  HS65_LL_NAND2X7 U11063 ( .A(n363), .B(n386), .Z(n7853) );
  HS65_LL_NAND2X7 U11064 ( .A(n165), .B(n149), .Z(n3572) );
  HS65_LL_NAND2X7 U11065 ( .A(n330), .B(n354), .Z(n8037) );
  HS65_LL_NAND2X7 U11066 ( .A(n653), .B(n635), .Z(n3334) );
  HS65_LL_NAND2X7 U11067 ( .A(n391), .B(n368), .Z(n8235) );
  HS65_LL_AOI12X2 U11068 ( .A(n77), .B(n59), .C(n6890), .Z(n6889) );
  HS65_LL_AOI12X2 U11069 ( .A(n259), .B(n236), .C(n5298), .Z(n5297) );
  HS65_LL_AOI12X2 U11070 ( .A(n301), .B(n278), .C(n7005), .Z(n7004) );
  HS65_LL_NAND2X7 U11071 ( .A(n345), .B(n328), .Z(n8348) );
  HS65_LL_NAND2X7 U11072 ( .A(n400), .B(n370), .Z(n8114) );
  HS65_LL_OAI21X3 U11073 ( .A(n851), .B(n845), .C(n875), .Z(n1438) );
  HS65_LL_OAI21X3 U11074 ( .A(n769), .B(n763), .C(n793), .Z(n2190) );
  HS65_LL_NAND2X7 U11075 ( .A(n341), .B(n335), .Z(n8537) );
  HS65_LL_NAND2X7 U11076 ( .A(n862), .B(n850), .Z(n1328) );
  HS65_LL_NAND2X7 U11077 ( .A(n780), .B(n768), .Z(n2080) );
  HS65_LL_AOI12X2 U11078 ( .A(n373), .B(n396), .C(n8284), .Z(n8283) );
  HS65_LL_NAND2X7 U11079 ( .A(n903), .B(n891), .Z(n2456) );
  HS65_LL_OAI21X3 U11080 ( .A(n892), .B(n886), .C(n916), .Z(n2566) );
  HS65_LL_NAND2X7 U11081 ( .A(n538), .B(n562), .Z(n6664) );
  HS65_LL_NAND2X7 U11082 ( .A(n16), .B(n40), .Z(n5071) );
  HS65_LL_NAND2X7 U11083 ( .A(n821), .B(n809), .Z(n1704) );
  HS65_LL_NAND2X7 U11084 ( .A(n246), .B(n255), .Z(n5281) );
  HS65_LL_NAND2X7 U11085 ( .A(n67), .B(n90), .Z(n6873) );
  HS65_LL_NAND2X7 U11086 ( .A(n377), .B(n386), .Z(n8262) );
  HS65_LL_OAI21X3 U11087 ( .A(n810), .B(n804), .C(n834), .Z(n1814) );
  HS65_LL_OAI21X3 U11088 ( .A(n914), .B(n906), .C(n891), .Z(n2571) );
  HS65_LL_NAND2X7 U11089 ( .A(n421), .B(n435), .Z(n3855) );
  HS65_LL_NAND2X7 U11090 ( .A(n190), .B(n223), .Z(n3500) );
  HS65_LL_OAI21X3 U11091 ( .A(n832), .B(n1594), .C(n802), .Z(n1628) );
  HS65_LL_OAI21X3 U11092 ( .A(n659), .B(n655), .C(n640), .Z(n4242) );
  HS65_LL_NAND2X7 U11093 ( .A(n396), .B(n368), .Z(n8289) );
  HS65_LL_NAND2X7 U11094 ( .A(n660), .B(n634), .Z(n3713) );
  HS65_LL_OAI21X3 U11095 ( .A(n914), .B(n2346), .C(n884), .Z(n2380) );
  HS65_LL_OAI21X3 U11096 ( .A(n873), .B(n1218), .C(n843), .Z(n1252) );
  HS65_LL_OAI21X3 U11097 ( .A(n791), .B(n1970), .C(n761), .Z(n2004) );
  HS65_LL_NAND2X7 U11098 ( .A(n793), .B(n768), .Z(n1902) );
  HS65_LL_NAND2X7 U11099 ( .A(n875), .B(n850), .Z(n1150) );
  HS65_LL_NAND2X7 U11100 ( .A(n639), .B(n648), .Z(n3740) );
  HS65_LL_OAI21X3 U11101 ( .A(n389), .B(n397), .C(n363), .Z(n8955) );
  HS65_LL_OAI21X3 U11102 ( .A(n349), .B(n343), .C(n323), .Z(n8863) );
  HS65_LL_NAND2X7 U11103 ( .A(n480), .B(n459), .Z(n5455) );
  HS65_LL_NAND2X7 U11104 ( .A(n263), .B(n242), .Z(n5340) );
  HS65_LL_NAND2X7 U11105 ( .A(n305), .B(n284), .Z(n7047) );
  HS65_LL_NAND2X7 U11106 ( .A(n86), .B(n54), .Z(n6932) );
  HS65_LL_NAND2X7 U11107 ( .A(n513), .B(n495), .Z(n6817) );
  HS65_LL_NAND2X7 U11108 ( .A(n689), .B(n671), .Z(n5225) );
  HS65_LL_NAND2X7 U11109 ( .A(n916), .B(n891), .Z(n2278) );
  HS65_LL_NAND2X7 U11110 ( .A(n834), .B(n809), .Z(n1526) );
  HS65_LL_OAI21X3 U11111 ( .A(n767), .B(n763), .C(n781), .Z(n2208) );
  HS65_LL_OAI21X3 U11112 ( .A(n849), .B(n845), .C(n863), .Z(n1456) );
  HS65_LL_NAND2X7 U11113 ( .A(n174), .B(n149), .Z(n3638) );
  HS65_LL_OAI21X3 U11114 ( .A(n890), .B(n886), .C(n904), .Z(n2584) );
  HS65_LL_NAND2X7 U11115 ( .A(n34), .B(n16), .Z(n5089) );
  HS65_LL_NAND2X7 U11116 ( .A(n556), .B(n538), .Z(n6682) );
  HS65_LL_NAND2X7 U11117 ( .A(n582), .B(n603), .Z(n8403) );
  HS65_LL_NAND2X7 U11118 ( .A(n102), .B(n123), .Z(n8455) );
  HS65_LL_OAI21X3 U11119 ( .A(n808), .B(n804), .C(n822), .Z(n1832) );
  HS65_LL_NAND2X7 U11120 ( .A(n422), .B(n435), .Z(n2999) );
  HS65_LL_NAND2X7 U11121 ( .A(n189), .B(n223), .Z(n2862) );
  HS65_LL_NAND2X7 U11122 ( .A(n356), .B(n335), .Z(n8591) );
  HS65_LL_IVX9 U11123 ( .A(n2821), .Z(n448) );
  HS65_LL_IVX9 U11124 ( .A(n2813), .Z(n273) );
  HS65_LL_NAND2X7 U11125 ( .A(n640), .B(n648), .Z(n2974) );
  HS65_LL_AOI12X2 U11126 ( .A(n770), .B(n787), .C(n2032), .Z(n2031) );
  HS65_LL_AOI12X2 U11127 ( .A(n852), .B(n869), .C(n1280), .Z(n1279) );
  HS65_LL_NAND2X7 U11128 ( .A(n172), .B(n151), .Z(n3600) );
  HS65_LL_AOI12X2 U11129 ( .A(n893), .B(n910), .C(n2408), .Z(n2407) );
  HS65_LL_NAND2X7 U11130 ( .A(n614), .B(n586), .Z(n8727) );
  HS65_LL_NAND2X7 U11131 ( .A(n134), .B(n106), .Z(n8817) );
  HS65_LL_NAND4ABX3 U11132 ( .A(n6065), .B(n6066), .C(n6067), .D(n6068), .Z(
        n6064) );
  HS65_LL_AOI212X4 U11133 ( .A(n537), .B(n555), .C(n532), .D(n569), .E(n6069), 
        .Z(n6068) );
  HS65_LL_NAND4ABX3 U11134 ( .A(n4472), .B(n4473), .C(n4474), .D(n4475), .Z(
        n4471) );
  HS65_LL_AOI212X4 U11135 ( .A(n15), .B(n33), .C(n10), .D(n47), .E(n4476), .Z(
        n4475) );
  HS65_LL_NAND4ABX3 U11136 ( .A(n4581), .B(n4582), .C(n4583), .D(n4584), .Z(
        n4580) );
  HS65_LL_AOI212X4 U11137 ( .A(n244), .B(n257), .C(n247), .D(n252), .E(n4585), 
        .Z(n4584) );
  HS65_LL_NAND4ABX3 U11138 ( .A(n6191), .B(n6192), .C(n6193), .D(n6194), .Z(
        n6190) );
  HS65_LL_AOI212X4 U11139 ( .A(n286), .B(n299), .C(n289), .D(n294), .E(n6195), 
        .Z(n6194) );
  HS65_LL_NAND4ABX3 U11140 ( .A(n6174), .B(n6175), .C(n6176), .D(n6177), .Z(
        n6173) );
  HS65_LL_AOI212X4 U11141 ( .A(n55), .B(n76), .C(n68), .D(n89), .E(n6178), .Z(
        n6177) );
  HS65_LL_NAND4ABX3 U11142 ( .A(n4598), .B(n4599), .C(n4600), .D(n4601), .Z(
        n4597) );
  HS65_LL_AOI212X4 U11143 ( .A(n461), .B(n474), .C(n464), .D(n469), .E(n4602), 
        .Z(n4601) );
  HS65_LL_NAND4ABX3 U11144 ( .A(n7998), .B(n7999), .C(n8000), .D(n8001), .Z(
        n7997) );
  HS65_LL_AOI212X4 U11145 ( .A(n614), .B(n578), .C(n583), .D(n602), .E(n8002), 
        .Z(n8001) );
  HS65_LL_NAND4ABX3 U11146 ( .A(n8011), .B(n8012), .C(n8013), .D(n8014), .Z(
        n8010) );
  HS65_LL_AOI212X4 U11147 ( .A(n134), .B(n98), .C(n103), .D(n122), .E(n8015), 
        .Z(n8014) );
  HS65_LL_NAND2X7 U11148 ( .A(n645), .B(n634), .Z(n3722) );
  HS65_LL_IVX9 U11149 ( .A(n7694), .Z(n575) );
  HS65_LL_NOR3AX2 U11150 ( .A(n7695), .B(n7696), .C(n7697), .Z(n7694) );
  HS65_LL_AO12X9 U11151 ( .A(n603), .B(n576), .C(n7698), .Z(n7696) );
  HS65_LL_IVX9 U11152 ( .A(n7732), .Z(n95) );
  HS65_LL_NOR3AX2 U11153 ( .A(n7733), .B(n7734), .C(n7735), .Z(n7732) );
  HS65_LL_AO12X9 U11154 ( .A(n123), .B(n96), .C(n7736), .Z(n7734) );
  HS65_LL_NAND2X7 U11155 ( .A(n600), .B(n591), .Z(n8718) );
  HS65_LL_NAND2X7 U11156 ( .A(n120), .B(n111), .Z(n8808) );
  HS65_LL_NOR4ABX2 U11157 ( .A(n6501), .B(n6479), .C(n6321), .D(n6178), .Z(
        n6828) );
  HS65_LL_NOR4ABX2 U11158 ( .A(n4908), .B(n4886), .C(n4741), .D(n4585), .Z(
        n5236) );
  HS65_LL_AOI12X2 U11159 ( .A(n654), .B(n634), .C(n3680), .Z(n3679) );
  HS65_LL_NAND2X7 U11160 ( .A(n244), .B(n260), .Z(n5280) );
  HS65_LL_NAND2X7 U11161 ( .A(n286), .B(n302), .Z(n6987) );
  HS65_LL_NAND2X7 U11162 ( .A(n55), .B(n83), .Z(n6872) );
  HS65_LL_NAND2X7 U11163 ( .A(n653), .B(n634), .Z(n3712) );
  HS65_LL_AOI12X2 U11164 ( .A(n63), .B(n90), .C(n6056), .Z(n6878) );
  HS65_LL_NOR4ABX2 U11165 ( .A(n2976), .B(n3144), .C(n3302), .D(n3312), .Z(
        n3656) );
  HS65_LL_NAND2X7 U11166 ( .A(n650), .B(n627), .Z(n3760) );
  HS65_LL_OAI21X3 U11167 ( .A(n842), .B(n1185), .C(n860), .Z(n1184) );
  HS65_LL_OAI21X3 U11168 ( .A(n760), .B(n1937), .C(n778), .Z(n1936) );
  HS65_LL_NAND2X7 U11169 ( .A(n441), .B(n408), .Z(n3875) );
  HS65_LL_NAND2X7 U11170 ( .A(n475), .B(n452), .Z(n4977) );
  HS65_LL_NAND2X7 U11171 ( .A(n258), .B(n235), .Z(n4924) );
  HS65_LL_NAND2X7 U11172 ( .A(n300), .B(n277), .Z(n6570) );
  HS65_LL_NAND2X7 U11173 ( .A(n73), .B(n66), .Z(n6517) );
  HS65_LL_NAND2X7 U11174 ( .A(n508), .B(n504), .Z(n6444) );
  HS65_LL_NAND2X7 U11175 ( .A(n684), .B(n680), .Z(n4851) );
  HS65_LL_NAND2X7 U11176 ( .A(n216), .B(n202), .Z(n2937) );
  HS65_LL_OAI21X3 U11177 ( .A(n883), .B(n2313), .C(n901), .Z(n2312) );
  HS65_LL_NAND2X7 U11178 ( .A(n814), .B(n828), .Z(n1675) );
  HS65_LL_NAND2X7 U11179 ( .A(n855), .B(n869), .Z(n1299) );
  HS65_LL_NAND2X7 U11180 ( .A(n773), .B(n787), .Z(n2051) );
  HS65_LL_NAND2X7 U11181 ( .A(n896), .B(n910), .Z(n2427) );
  HS65_LL_OAI21X3 U11182 ( .A(n801), .B(n1561), .C(n819), .Z(n1560) );
  HS65_LL_NAND2X7 U11183 ( .A(n429), .B(n416), .Z(n3828) );
  HS65_LL_NAND2X7 U11184 ( .A(n210), .B(n195), .Z(n3472) );
  HS65_LL_NAND2X7 U11185 ( .A(n37), .B(n25), .Z(n5096) );
  HS65_LL_NAND2X7 U11186 ( .A(n559), .B(n547), .Z(n6689) );
  HS65_LL_NOR4ABX2 U11187 ( .A(n8069), .B(n7862), .C(n8093), .D(n7974), .Z(
        n8191) );
  HS65_LL_NAND2X7 U11188 ( .A(n659), .B(n627), .Z(n3759) );
  HS65_LL_NAND2X7 U11189 ( .A(n29), .B(n25), .Z(n4713) );
  HS65_LL_NAND2X7 U11190 ( .A(n551), .B(n547), .Z(n6306) );
  HS65_LL_NOR4ABX2 U11191 ( .A(n7771), .B(n7772), .C(n7773), .D(n7774), .Z(
        n7757) );
  HS65_LL_NOR4ABX2 U11192 ( .A(n7101), .B(n7236), .C(n7237), .D(n7067), .Z(
        n7230) );
  HS65_LL_IVX9 U11193 ( .A(n2783), .Z(n51) );
  HS65_LL_IVX9 U11194 ( .A(n2791), .Z(n229) );
  HS65_LL_NAND2X7 U11195 ( .A(n436), .B(n408), .Z(n3202) );
  HS65_LL_NAND2X7 U11196 ( .A(n391), .B(n376), .Z(n8300) );
  HS65_LL_NOR4ABX2 U11197 ( .A(n7753), .B(n7754), .C(n7755), .D(n7756), .Z(
        n7739) );
  HS65_LL_NOR3AX2 U11198 ( .A(n2975), .B(n3302), .C(n3145), .Z(n3287) );
  HS65_LL_NOR4ABX2 U11199 ( .A(n3946), .B(n3947), .C(n3948), .D(n3949), .Z(
        n3942) );
  HS65_LL_MX41X7 U11200 ( .D0(n660), .S0(n633), .D1(n627), .S1(n655), .D2(n652), .S2(n631), .D3(n629), .S3(n644), .Z(n3949) );
  HS65_LL_NOR4ABX2 U11201 ( .A(n3966), .B(n3967), .C(n3968), .D(n3969), .Z(
        n3962) );
  HS65_LL_MX41X7 U11202 ( .D0(n429), .S0(n415), .D1(n408), .S1(n438), .D2(n443), .S2(n413), .D3(n411), .S3(n431), .Z(n3969) );
  HS65_LL_NAND2X7 U11203 ( .A(n640), .B(n658), .Z(n3726) );
  HS65_LL_NAND2X7 U11204 ( .A(n428), .B(n408), .Z(n3874) );
  HS65_LL_NAND2X7 U11205 ( .A(n814), .B(n829), .Z(n1740) );
  HS65_LL_NOR4ABX2 U11206 ( .A(n7184), .B(n7120), .C(n6044), .D(n7115), .Z(
        n7411) );
  HS65_LL_NAND2X7 U11207 ( .A(n773), .B(n788), .Z(n2116) );
  HS65_LL_NAND2X7 U11208 ( .A(n855), .B(n870), .Z(n1364) );
  HS65_LL_NAND2X7 U11209 ( .A(n896), .B(n911), .Z(n2492) );
  HS65_LL_NAND2X7 U11210 ( .A(n220), .B(n196), .Z(n3529) );
  HS65_LL_NAND2X7 U11211 ( .A(n371), .B(n384), .Z(n8239) );
  HS65_LL_NAND2X7 U11212 ( .A(n324), .B(n345), .Z(n8541) );
  HS65_LL_NAND2X7 U11213 ( .A(n429), .B(n412), .Z(n3804) );
  HS65_LL_NAND2X7 U11214 ( .A(n210), .B(n199), .Z(n3447) );
  HS65_LL_NAND2X7 U11215 ( .A(n343), .B(n327), .Z(n8608) );
  HS65_LL_NAND2X7 U11216 ( .A(n871), .B(n839), .Z(n1303) );
  HS65_LL_NAND2X7 U11217 ( .A(n789), .B(n757), .Z(n2055) );
  HS65_LL_NAND2X7 U11218 ( .A(n267), .B(n241), .Z(n4752) );
  HS65_LL_NAND2X7 U11219 ( .A(n520), .B(n493), .Z(n6226) );
  HS65_LL_NAND2X7 U11220 ( .A(n484), .B(n458), .Z(n4779) );
  HS65_LL_NAND2X7 U11221 ( .A(n309), .B(n283), .Z(n6372) );
  HS65_LL_NAND2X7 U11222 ( .A(n81), .B(n57), .Z(n6333) );
  HS65_LL_NAND2X7 U11223 ( .A(n696), .B(n669), .Z(n4633) );
  HS65_LL_NOR3AX2 U11224 ( .A(n2848), .B(n2849), .C(n2850), .Z(n2825) );
  HS65_LL_NAND2X7 U11225 ( .A(n848), .B(n869), .Z(n1298) );
  HS65_LL_NAND2X7 U11226 ( .A(n766), .B(n787), .Z(n2050) );
  HS65_LL_NAND2X7 U11227 ( .A(n261), .B(n241), .Z(n4931) );
  HS65_LL_NAND2X7 U11228 ( .A(n478), .B(n458), .Z(n4984) );
  HS65_LL_NAND2X7 U11229 ( .A(n303), .B(n283), .Z(n6577) );
  HS65_LL_NAND2X7 U11230 ( .A(n85), .B(n57), .Z(n6524) );
  HS65_LL_NAND2X7 U11231 ( .A(n516), .B(n493), .Z(n6451) );
  HS65_LL_NAND2X7 U11232 ( .A(n692), .B(n669), .Z(n4858) );
  HS65_LL_NAND2X7 U11233 ( .A(n31), .B(n22), .Z(n5065) );
  HS65_LL_NAND2X7 U11234 ( .A(n553), .B(n544), .Z(n6658) );
  HS65_LL_NAND2X7 U11235 ( .A(n363), .B(n390), .Z(n8249) );
  HS65_LL_NAND2X7 U11236 ( .A(n830), .B(n798), .Z(n1679) );
  HS65_LL_NAND2X7 U11237 ( .A(n912), .B(n880), .Z(n2431) );
  HS65_LL_NAND2X7 U11238 ( .A(n889), .B(n910), .Z(n2426) );
  HS65_LL_NAND2X7 U11239 ( .A(n660), .B(n630), .Z(n3689) );
  HS65_LL_NAND2X7 U11240 ( .A(n371), .B(n400), .Z(n8246) );
  HS65_LL_AOI12X2 U11241 ( .A(n245), .B(n4927), .C(n4928), .Z(n4926) );
  HS65_LL_AOI12X2 U11242 ( .A(n69), .B(n6520), .C(n6521), .Z(n6519) );
  HS65_LL_NAND2X7 U11243 ( .A(n216), .B(n195), .Z(n3471) );
  HS65_LL_NAND2X7 U11244 ( .A(n807), .B(n828), .Z(n1674) );
  HS65_LL_NAND2X7 U11245 ( .A(n649), .B(n628), .Z(n3768) );
  HS65_LL_NAND2X7 U11246 ( .A(n905), .B(n890), .Z(n2451) );
  HS65_LL_NAND2X7 U11247 ( .A(n864), .B(n849), .Z(n1323) );
  HS65_LL_NAND2X7 U11248 ( .A(n782), .B(n767), .Z(n2075) );
  HS65_LL_NAND2X7 U11249 ( .A(n823), .B(n808), .Z(n1699) );
  HS65_LL_NAND2X7 U11250 ( .A(n419), .B(n440), .Z(n3850) );
  HS65_LL_NOR3AX2 U11251 ( .A(n4672), .B(n4544), .C(n4473), .Z(n4655) );
  HS65_LL_NOR3AX2 U11252 ( .A(n6265), .B(n6137), .C(n6066), .Z(n6248) );
  HS65_LL_NOR3AX2 U11253 ( .A(n6479), .B(n6322), .C(n6175), .Z(n6463) );
  HS65_LL_NOR3AX2 U11254 ( .A(n4886), .B(n4742), .C(n4582), .Z(n4870) );
  HS65_LL_NAND2X7 U11255 ( .A(n637), .B(n649), .Z(n3735) );
  HS65_LL_NAND2X7 U11256 ( .A(n436), .B(n416), .Z(n3827) );
  HS65_LL_OAI21X3 U11257 ( .A(n340), .B(n352), .C(n320), .Z(n8895) );
  HS65_LL_NAND2X7 U11258 ( .A(n823), .B(n798), .Z(n1605) );
  HS65_LL_NAND2X7 U11259 ( .A(n782), .B(n757), .Z(n1981) );
  HS65_LL_NAND2X7 U11260 ( .A(n864), .B(n839), .Z(n1229) );
  HS65_LL_NAND2X7 U11261 ( .A(n905), .B(n880), .Z(n2357) );
  HS65_LL_NOR4ABX2 U11262 ( .A(n3029), .B(n3638), .C(n3274), .D(n3246), .Z(
        n4141) );
  HS65_LL_OAI21X3 U11263 ( .A(n580), .B(n579), .C(n599), .Z(n7795) );
  HS65_LL_OAI21X3 U11264 ( .A(n100), .B(n99), .C(n119), .Z(n7894) );
  HS65_LL_OAI21X3 U11265 ( .A(n635), .B(n633), .C(n648), .Z(n4247) );
  HS65_LL_NOR4ABX2 U11266 ( .A(n3652), .B(n3653), .C(n3654), .D(n3655), .Z(
        n3640) );
  HS65_LL_NAND2X7 U11267 ( .A(n538), .B(n557), .Z(n6665) );
  HS65_LL_NAND2X7 U11268 ( .A(n16), .B(n35), .Z(n5072) );
  HS65_LL_NAND2X7 U11269 ( .A(n111), .B(n127), .Z(n8774) );
  HS65_LL_NAND2X7 U11270 ( .A(n591), .B(n607), .Z(n8684) );
  HS65_LL_NAND2X7 U11271 ( .A(n576), .B(n617), .Z(n8699) );
  HS65_LL_NOR3AX2 U11272 ( .A(n2337), .B(n2348), .C(n2302), .Z(n2420) );
  HS65_LL_NOR3AX2 U11273 ( .A(n1209), .B(n1220), .C(n1174), .Z(n1292) );
  HS65_LL_NOR3AX2 U11274 ( .A(n1961), .B(n1972), .C(n1926), .Z(n2044) );
  HS65_LL_NOR3AX2 U11275 ( .A(n1585), .B(n1596), .C(n1550), .Z(n1668) );
  HS65_LL_NOR3AX2 U11276 ( .A(n3355), .B(n3367), .C(n3169), .Z(n3821) );
  HS65_LL_NOR3AX2 U11277 ( .A(n3070), .B(n3082), .C(n2942), .Z(n3465) );
  HS65_LL_NOR4ABX2 U11278 ( .A(n1764), .B(n1765), .C(n1766), .D(n1767), .Z(
        n1760) );
  HS65_LL_MX41X7 U11279 ( .D0(n814), .S0(n824), .D1(n826), .S1(n804), .D2(n799), .S2(n825), .D3(n831), .S3(n802), .Z(n1767) );
  HS65_LL_NOR4ABX2 U11280 ( .A(n2140), .B(n2141), .C(n2142), .D(n2143), .Z(
        n2136) );
  HS65_LL_MX41X7 U11281 ( .D0(n773), .S0(n783), .D1(n785), .S1(n763), .D2(n758), .S2(n784), .D3(n790), .S3(n761), .Z(n2143) );
  HS65_LL_NOR4ABX2 U11282 ( .A(n1388), .B(n1389), .C(n1390), .D(n1391), .Z(
        n1384) );
  HS65_LL_MX41X7 U11283 ( .D0(n855), .S0(n865), .D1(n867), .S1(n845), .D2(n840), .S2(n866), .D3(n872), .S3(n843), .Z(n1391) );
  HS65_LL_NOR4ABX2 U11284 ( .A(n2516), .B(n2517), .C(n2518), .D(n2519), .Z(
        n2512) );
  HS65_LL_MX41X7 U11285 ( .D0(n896), .S0(n906), .D1(n908), .S1(n886), .D2(n881), .S2(n907), .D3(n913), .S3(n884), .Z(n2519) );
  HS65_LL_NOR4ABX2 U11286 ( .A(n4064), .B(n4050), .C(n3921), .D(n4191), .Z(
        n4187) );
  HS65_LL_MX41X7 U11287 ( .D0(n210), .S0(n192), .D1(n202), .S1(n214), .D2(n218), .S2(n198), .D3(n197), .S3(n225), .Z(n4191) );
  HS65_LL_NOR4ABX2 U11288 ( .A(n1919), .B(n2090), .C(n1954), .D(n2015), .Z(
        n2199) );
  HS65_LL_NOR4ABX2 U11289 ( .A(n1167), .B(n1338), .C(n1202), .D(n1263), .Z(
        n1447) );
  HS65_LL_OAI21X3 U11290 ( .A(n370), .B(n367), .C(n386), .Z(n8960) );
  HS65_LL_NOR4ABX2 U11291 ( .A(n2863), .B(n2864), .C(n2865), .D(n2866), .Z(
        n2852) );
  HS65_LL_AO212X4 U11292 ( .A(n193), .B(n221), .C(n189), .D(n226), .E(n2867), 
        .Z(n2865) );
  HS65_LL_NAND2X7 U11293 ( .A(n386), .B(n365), .Z(n8263) );
  HS65_LL_NAND2X7 U11294 ( .A(n347), .B(n319), .Z(n8565) );
  HS65_LL_NOR4ABX2 U11295 ( .A(n2975), .B(n2976), .C(n2977), .D(n2978), .Z(
        n2965) );
  HS65_LL_AO212X4 U11296 ( .A(n636), .B(n650), .C(n640), .D(n645), .E(n2979), 
        .Z(n2977) );
  HS65_LL_NOR4ABX2 U11297 ( .A(n5096), .B(n5097), .C(n5098), .D(n5099), .Z(
        n5084) );
  HS65_LL_NOR4ABX2 U11298 ( .A(n6689), .B(n6690), .C(n6691), .D(n6692), .Z(
        n6677) );
  HS65_LL_NOR4ABX2 U11299 ( .A(n1543), .B(n1714), .C(n1578), .D(n1639), .Z(
        n1823) );
  HS65_LL_NOR4ABX2 U11300 ( .A(n2295), .B(n2466), .C(n2330), .D(n2391), .Z(
        n2575) );
  HS65_LL_NOR3AX2 U11301 ( .A(n7249), .B(n7250), .C(n7069), .Z(n7243) );
  HS65_LL_AO12X9 U11302 ( .A(n568), .B(n538), .C(n7256), .Z(n7250) );
  HS65_LL_NOR3AX2 U11303 ( .A(n5657), .B(n5658), .C(n5477), .Z(n5651) );
  HS65_LL_AO12X9 U11304 ( .A(n46), .B(n16), .C(n5664), .Z(n5658) );
  HS65_LL_NOR3AX2 U11305 ( .A(n4510), .B(n5905), .C(n5557), .Z(n5899) );
  HS65_LL_AO12X9 U11306 ( .A(n467), .B(n459), .C(n5553), .Z(n5905) );
  HS65_LL_NOR3AX2 U11307 ( .A(n6103), .B(n7497), .C(n7149), .Z(n7491) );
  HS65_LL_AO12X9 U11308 ( .A(n292), .B(n284), .C(n7145), .Z(n7497) );
  HS65_LL_NOR3AX2 U11309 ( .A(n4449), .B(n5846), .C(n5535), .Z(n5840) );
  HS65_LL_AO12X9 U11310 ( .A(n250), .B(n242), .C(n5531), .Z(n5846) );
  HS65_LL_NOR3AX2 U11311 ( .A(n6042), .B(n7438), .C(n7127), .Z(n7432) );
  HS65_LL_AO12X9 U11312 ( .A(n91), .B(n54), .C(n7123), .Z(n7438) );
  HS65_LL_NOR3AX2 U11313 ( .A(n5687), .B(n5688), .C(n5491), .Z(n5681) );
  HS65_LL_AO12X9 U11314 ( .A(n701), .B(n671), .C(n5694), .Z(n5688) );
  HS65_LL_NOR3AX2 U11315 ( .A(n7279), .B(n7280), .C(n7083), .Z(n7273) );
  HS65_LL_AO12X9 U11316 ( .A(n525), .B(n495), .C(n7286), .Z(n7280) );
  HS65_LL_OAI21X3 U11317 ( .A(n334), .B(n333), .C(n347), .Z(n8900) );
  HS65_LL_NOR4ABX2 U11318 ( .A(n2450), .B(n2332), .C(n2478), .D(n2461), .Z(
        n2543) );
  HS65_LL_NOR4ABX2 U11319 ( .A(n8591), .B(n8592), .C(n8593), .D(n8594), .Z(
        n8579) );
  HS65_LL_NAND2X7 U11320 ( .A(n495), .B(n514), .Z(n6785) );
  HS65_LL_NAND2X7 U11321 ( .A(n671), .B(n690), .Z(n5193) );
  HS65_LL_NAND2X7 U11322 ( .A(n54), .B(n83), .Z(n6901) );
  HS65_LL_NAND2X7 U11323 ( .A(n242), .B(n260), .Z(n5309) );
  HS65_LL_NAND2X7 U11324 ( .A(n459), .B(n477), .Z(n5424) );
  HS65_LL_NAND2X7 U11325 ( .A(n284), .B(n302), .Z(n7016) );
  HS65_LL_NOR4ABX2 U11326 ( .A(n2074), .B(n1956), .C(n2102), .D(n2085), .Z(
        n2167) );
  HS65_LL_NOR4ABX2 U11327 ( .A(n5415), .B(n5424), .C(n5393), .D(n4969), .Z(
        n5926) );
  HS65_LL_NOR4ABX2 U11328 ( .A(n7007), .B(n7016), .C(n6985), .D(n6562), .Z(
        n7518) );
  HS65_LL_NOR4ABX2 U11329 ( .A(n5300), .B(n5309), .C(n5278), .D(n4916), .Z(
        n5867) );
  HS65_LL_NOR4ABX2 U11330 ( .A(n6892), .B(n6901), .C(n6870), .D(n6509), .Z(
        n7463) );
  HS65_LL_NOR4ABX2 U11331 ( .A(n5184), .B(n5193), .C(n5161), .D(n4841), .Z(
        n5763) );
  HS65_LL_NOR4ABX2 U11332 ( .A(n6776), .B(n6785), .C(n6753), .D(n6434), .Z(
        n7355) );
  HS65_LL_NOR4ABX2 U11333 ( .A(n1698), .B(n1580), .C(n1726), .D(n1709), .Z(
        n1791) );
  HS65_LL_NOR4ABX2 U11334 ( .A(n5405), .B(n5455), .C(n4960), .D(n4947), .Z(
        n5626) );
  HS65_LL_NOR4ABX2 U11335 ( .A(n5290), .B(n5340), .C(n4907), .D(n4894), .Z(
        n5601) );
  HS65_LL_NOR4ABX2 U11336 ( .A(n6997), .B(n7047), .C(n6553), .D(n6540), .Z(
        n7218) );
  HS65_LL_NOR4ABX2 U11337 ( .A(n5174), .B(n5225), .C(n4832), .D(n4819), .Z(
        n5792) );
  HS65_LL_NOR4ABX2 U11338 ( .A(n6766), .B(n6817), .C(n6425), .D(n6412), .Z(
        n7384) );
  HS65_LL_NOR4ABX2 U11339 ( .A(n6882), .B(n6932), .C(n6500), .D(n6487), .Z(
        n7193) );
  HS65_LL_NAND2X7 U11340 ( .A(n350), .B(n322), .Z(n8514) );
  HS65_LL_NOR4ABX2 U11341 ( .A(n8289), .B(n8290), .C(n8291), .D(n8292), .Z(
        n8277) );
  HS65_LL_NOR4ABX2 U11342 ( .A(n8114), .B(n8074), .C(n8265), .D(n8223), .Z(
        n8981) );
  HS65_LL_NOR4ABX2 U11343 ( .A(n3734), .B(n3298), .C(n3762), .D(n3745), .Z(
        n4015) );
  HS65_LL_NOR4ABX2 U11344 ( .A(n8711), .B(n7796), .C(n7690), .D(n8712), .Z(
        n8705) );
  HS65_LL_NOR4ABX2 U11345 ( .A(n8801), .B(n7895), .C(n7728), .D(n8802), .Z(
        n8795) );
  HS65_LL_NOR4ABX2 U11346 ( .A(n5343), .B(n5344), .C(n5345), .D(n5346), .Z(
        n5336) );
  HS65_LL_NOR4ABX2 U11347 ( .A(n5458), .B(n5459), .C(n5460), .D(n5461), .Z(
        n5451) );
  HS65_LL_NOR4ABX2 U11348 ( .A(n7050), .B(n7051), .C(n7052), .D(n7053), .Z(
        n7043) );
  HS65_LL_NOR4ABX2 U11349 ( .A(n6935), .B(n6936), .C(n6937), .D(n6938), .Z(
        n6928) );
  HS65_LL_NOR4ABX2 U11350 ( .A(n3763), .B(n3764), .C(n3765), .D(n3766), .Z(
        n3756) );
  HS65_LL_NOR4ABX2 U11351 ( .A(n2595), .B(n2480), .C(n2368), .D(n2399), .Z(
        n2589) );
  HS65_LL_OAI21X3 U11352 ( .A(n904), .B(n905), .C(n895), .Z(n2595) );
  HS65_LL_NOR4ABX2 U11353 ( .A(n1731), .B(n1732), .C(n1733), .D(n1734), .Z(
        n1719) );
  HS65_LL_NOR4ABX2 U11354 ( .A(n1186), .B(n1187), .C(n1188), .D(n1189), .Z(
        n1176) );
  HS65_LL_NOR4ABX2 U11355 ( .A(n1938), .B(n1939), .C(n1940), .D(n1941), .Z(
        n1928) );
  HS65_LL_NOR4ABX2 U11356 ( .A(n2219), .B(n2104), .C(n1992), .D(n2023), .Z(
        n2213) );
  HS65_LL_OAI21X3 U11357 ( .A(n781), .B(n782), .C(n772), .Z(n2219) );
  HS65_LL_NOR4ABX2 U11358 ( .A(n1467), .B(n1352), .C(n1240), .D(n1271), .Z(
        n1461) );
  HS65_LL_OAI21X3 U11359 ( .A(n863), .B(n864), .C(n854), .Z(n1467) );
  HS65_LL_NOR4ABX2 U11360 ( .A(n2483), .B(n2484), .C(n2485), .D(n2486), .Z(
        n2471) );
  HS65_LL_NOR4ABX2 U11361 ( .A(n2314), .B(n2315), .C(n2316), .D(n2317), .Z(
        n2304) );
  HS65_LL_NOR4ABX2 U11362 ( .A(n1355), .B(n1356), .C(n1357), .D(n1358), .Z(
        n1343) );
  HS65_LL_NOR4ABX2 U11363 ( .A(n2107), .B(n2108), .C(n2109), .D(n2110), .Z(
        n2095) );
  HS65_LL_NAND2X7 U11364 ( .A(n399), .B(n366), .Z(n8211) );
  HS65_LL_NOR4ABX2 U11365 ( .A(n3882), .B(n3883), .C(n3884), .D(n3885), .Z(
        n3870) );
  HS65_LL_NOR4ABX2 U11366 ( .A(n6518), .B(n6474), .C(n6860), .D(n6880), .Z(
        n7198) );
  HS65_LL_NOR4ABX2 U11367 ( .A(n8454), .B(n8786), .C(n8820), .D(n8464), .Z(
        n9074) );
  HS65_LL_NOR4ABX2 U11368 ( .A(n8402), .B(n8696), .C(n8730), .D(n8412), .Z(
        n9016) );
  HS65_LL_NOR4ABX2 U11369 ( .A(n4200), .B(n3525), .C(n3104), .D(n3428), .Z(
        n4197) );
  HS65_LL_OAI21X3 U11370 ( .A(n193), .B(n191), .C(n219), .Z(n4200) );
  HS65_LL_NOR4ABX2 U11371 ( .A(n6654), .B(n6655), .C(n6656), .D(n6657), .Z(
        n6647) );
  HS65_LL_NOR4ABX2 U11372 ( .A(n5061), .B(n5062), .C(n5063), .D(n5064), .Z(
        n5054) );
  HS65_LL_NOR4ABX2 U11373 ( .A(n3689), .B(n3151), .C(n3711), .D(n3320), .Z(
        n4010) );
  HS65_LL_NOR4ABX2 U11374 ( .A(n3528), .B(n3471), .C(n3509), .D(n3094), .Z(
        n4170) );
  HS65_LL_OAI21X3 U11375 ( .A(n759), .B(n760), .C(n778), .Z(n2139) );
  HS65_LL_NOR3AX2 U11376 ( .A(n1566), .B(n1567), .C(n1568), .Z(n1551) );
  HS65_LL_NOR4ABX2 U11377 ( .A(n8290), .B(n8267), .C(n8232), .D(n8105), .Z(
        n8957) );
  HS65_LL_OAI21X3 U11378 ( .A(n841), .B(n842), .C(n860), .Z(n1387) );
  HS65_LL_OAI21X3 U11379 ( .A(n800), .B(n801), .C(n819), .Z(n1763) );
  HS65_LL_OAI21X3 U11380 ( .A(n882), .B(n883), .C(n901), .Z(n2515) );
  HS65_LL_NOR4ABX2 U11381 ( .A(n8239), .B(n8282), .C(n8206), .D(n8274), .Z(
        n8952) );
  HS65_LL_NOR4ABX2 U11382 ( .A(n3528), .B(n3529), .C(n3530), .D(n3531), .Z(
        n3516) );
  HS65_LL_NOR4ABX2 U11383 ( .A(n6775), .B(n6776), .C(n6777), .D(n6778), .Z(
        n6768) );
  HS65_LL_NOR4ABX2 U11384 ( .A(n5183), .B(n5184), .C(n5185), .D(n5186), .Z(
        n5176) );
  HS65_LL_NOR4ABX2 U11385 ( .A(n6891), .B(n6892), .C(n6893), .D(n6894), .Z(
        n6884) );
  HS65_LL_NOR4ABX2 U11386 ( .A(n5299), .B(n5300), .C(n5301), .D(n5302), .Z(
        n5292) );
  HS65_LL_NOR4ABX2 U11387 ( .A(n5414), .B(n5415), .C(n5416), .D(n5417), .Z(
        n5407) );
  HS65_LL_NOR4ABX2 U11388 ( .A(n7006), .B(n7007), .C(n7008), .D(n7009), .Z(
        n6999) );
  HS65_LL_NOR4ABX2 U11389 ( .A(n8592), .B(n8336), .C(n8534), .D(n8571), .Z(
        n8897) );
  HS65_LL_NAND2X7 U11390 ( .A(n792), .B(n759), .Z(n1977) );
  HS65_LL_NAND2X7 U11391 ( .A(n874), .B(n841), .Z(n1225) );
  HS65_LL_NAND2X7 U11392 ( .A(n833), .B(n800), .Z(n1601) );
  HS65_LL_NAND2X7 U11393 ( .A(n915), .B(n882), .Z(n2353) );
  HS65_LL_NOR4ABX2 U11394 ( .A(n2937), .B(n3511), .C(n3064), .D(n3419), .Z(
        n4207) );
  HS65_LL_NOR4ABX2 U11395 ( .A(n3202), .B(n3865), .C(n3409), .D(n3778), .Z(
        n4310) );
  HS65_LL_NAND2X7 U11396 ( .A(n282), .B(n299), .Z(n7006) );
  HS65_LL_NAND2X7 U11397 ( .A(n62), .B(n76), .Z(n6891) );
  HS65_LL_NAND2X7 U11398 ( .A(n240), .B(n257), .Z(n5299) );
  HS65_LL_NAND2X7 U11399 ( .A(n457), .B(n474), .Z(n5414) );
  HS65_LL_NOR4ABX2 U11400 ( .A(n8541), .B(n8584), .C(n8509), .D(n8575), .Z(
        n8892) );
  HS65_LL_NAND2X7 U11401 ( .A(n543), .B(n555), .Z(n6655) );
  HS65_LL_NAND2X7 U11402 ( .A(n21), .B(n33), .Z(n5062) );
  HS65_LL_NOR4ABX2 U11403 ( .A(n8347), .B(n8359), .C(n8567), .D(n8600), .Z(
        n8913) );
  HS65_LL_NOR3AX2 U11404 ( .A(n3347), .B(n3348), .C(n3349), .Z(n3336) );
  HS65_LL_OAI21X3 U11405 ( .A(n635), .B(n3311), .C(n644), .Z(n3347) );
  HS65_LL_NOR4ABX2 U11406 ( .A(n7796), .B(n7797), .C(n7798), .D(n7799), .Z(
        n7785) );
  HS65_LL_NOR4ABX2 U11407 ( .A(n7895), .B(n7896), .C(n7897), .D(n7898), .Z(
        n7884) );
  HS65_LL_NAND2X7 U11408 ( .A(n110), .B(n130), .Z(n8803) );
  HS65_LL_NAND2X7 U11409 ( .A(n590), .B(n610), .Z(n8713) );
  HS65_LL_NOR4ABX2 U11410 ( .A(n6654), .B(n6665), .C(n6633), .D(n6296), .Z(
        n7293) );
  HS65_LL_NOR4ABX2 U11411 ( .A(n5061), .B(n5072), .C(n5040), .D(n4703), .Z(
        n5701) );
  HS65_LL_NAND2X7 U11412 ( .A(n369), .B(n400), .Z(n8266) );
  HS65_LL_NOR4ABX2 U11413 ( .A(n3389), .B(n3856), .C(n3787), .D(n3400), .Z(
        n4034) );
  HS65_LL_NOR4ABX2 U11414 ( .A(n8862), .B(n8348), .C(n8590), .D(n8599), .Z(
        n8859) );
  HS65_LL_OAI21X3 U11415 ( .A(n332), .B(n317), .C(n356), .Z(n8862) );
  HS65_LL_NAND2X7 U11416 ( .A(n245), .B(n261), .Z(n5320) );
  HS65_LL_NAND2X7 U11417 ( .A(n462), .B(n478), .Z(n5435) );
  HS65_LL_NAND2X7 U11418 ( .A(n69), .B(n85), .Z(n6912) );
  HS65_LL_NAND2X7 U11419 ( .A(n287), .B(n303), .Z(n7027) );
  HS65_LL_NAND4ABX3 U11420 ( .A(n3296), .B(n3662), .C(n3139), .D(n3750), .Z(
        n4251) );
  HS65_LL_NAND4ABX3 U11421 ( .A(n1546), .B(n1547), .C(n1513), .D(n1548), .Z(
        n1528) );
  HS65_LL_AOI212X4 U11422 ( .A(n827), .B(n800), .C(n824), .D(n813), .E(n1549), 
        .Z(n1548) );
  HS65_LL_AO12X9 U11423 ( .A(n819), .B(n799), .C(n1550), .Z(n1549) );
  HS65_LL_NAND4ABX3 U11424 ( .A(n1922), .B(n1923), .C(n1889), .D(n1924), .Z(
        n1904) );
  HS65_LL_AOI212X4 U11425 ( .A(n786), .B(n759), .C(n783), .D(n772), .E(n1925), 
        .Z(n1924) );
  HS65_LL_AO12X9 U11426 ( .A(n778), .B(n758), .C(n1926), .Z(n1925) );
  HS65_LL_NAND4ABX3 U11427 ( .A(n1170), .B(n1171), .C(n1137), .D(n1172), .Z(
        n1152) );
  HS65_LL_AOI212X4 U11428 ( .A(n868), .B(n841), .C(n865), .D(n854), .E(n1173), 
        .Z(n1172) );
  HS65_LL_AO12X9 U11429 ( .A(n860), .B(n840), .C(n1174), .Z(n1173) );
  HS65_LL_NAND4ABX3 U11430 ( .A(n2298), .B(n2299), .C(n2265), .D(n2300), .Z(
        n2280) );
  HS65_LL_AOI212X4 U11431 ( .A(n909), .B(n882), .C(n906), .D(n895), .E(n2301), 
        .Z(n2300) );
  HS65_LL_AO12X9 U11432 ( .A(n901), .B(n881), .C(n2302), .Z(n2301) );
  HS65_LL_NOR4ABX2 U11433 ( .A(n4139), .B(n3572), .C(n3557), .D(n3582), .Z(
        n4134) );
  HS65_LL_OAI21X3 U11434 ( .A(n148), .B(n146), .C(n164), .Z(n4139) );
  HS65_LL_NAND4ABX3 U11435 ( .A(n8120), .B(n8268), .C(n8197), .D(n7970), .Z(
        n8949) );
  HS65_LL_NOR4ABX2 U11436 ( .A(n5052), .B(n5089), .C(n4694), .D(n4680), .Z(
        n5730) );
  HS65_LL_NOR4ABX2 U11437 ( .A(n6645), .B(n6682), .C(n6287), .D(n6273), .Z(
        n7322) );
  HS65_LL_NAND2X7 U11438 ( .A(n384), .B(n376), .Z(n8115) );
  HS65_LL_NAND2X7 U11439 ( .A(n855), .B(n871), .Z(n1355) );
  HS65_LL_NAND2X7 U11440 ( .A(n773), .B(n789), .Z(n2107) );
  HS65_LL_NAND2X7 U11441 ( .A(n429), .B(n407), .Z(n3882) );
  HS65_LLS_XOR3X2 U11442 ( .A(n2666), .B(n2628), .C(n2702), .Z(n2737) );
  HS65_LL_NAND2X7 U11443 ( .A(n371), .B(n391), .Z(n8290) );
  HS65_LL_NAND2X7 U11444 ( .A(n896), .B(n912), .Z(n2483) );
  HS65_LL_NAND2X7 U11445 ( .A(n814), .B(n830), .Z(n1731) );
  HS65_LL_NAND2X7 U11446 ( .A(n480), .B(n460), .Z(n5418) );
  HS65_LL_NAND2X7 U11447 ( .A(n263), .B(n243), .Z(n5303) );
  HS65_LL_NAND2X7 U11448 ( .A(n305), .B(n285), .Z(n7010) );
  HS65_LL_NAND2X7 U11449 ( .A(n689), .B(n672), .Z(n5187) );
  HS65_LL_NAND2X7 U11450 ( .A(n513), .B(n496), .Z(n6779) );
  HS65_LL_NAND2X7 U11451 ( .A(n86), .B(n56), .Z(n6895) );
  HS65_LL_NAND2X7 U11452 ( .A(n210), .B(n200), .Z(n3528) );
  HS65_LL_NAND2X7 U11453 ( .A(n324), .B(n341), .Z(n8592) );
  HS65_LL_NAND2X7 U11454 ( .A(n660), .B(n626), .Z(n3767) );
  HS65_LL_NAND2X7 U11455 ( .A(n913), .B(n890), .Z(n2315) );
  HS65_LL_NAND2X7 U11456 ( .A(n790), .B(n767), .Z(n1939) );
  HS65_LL_NAND2X7 U11457 ( .A(n872), .B(n849), .Z(n1187) );
  HS65_LL_NAND2X7 U11458 ( .A(n831), .B(n808), .Z(n1563) );
  HS65_LL_NAND2X7 U11459 ( .A(n411), .B(n440), .Z(n3177) );
  HS65_LL_NAND2X7 U11460 ( .A(n197), .B(n220), .Z(n2950) );
  HS65_LL_NAND2X7 U11461 ( .A(n180), .B(n155), .Z(n3653) );
  HS65_LL_NAND2X7 U11462 ( .A(n907), .B(n889), .Z(n2480) );
  HS65_LL_NAND2X7 U11463 ( .A(n629), .B(n649), .Z(n3151) );
  HS65_LL_NAND2X7 U11464 ( .A(n155), .B(n173), .Z(n3652) );
  HS65_LL_NAND2X7 U11465 ( .A(n451), .B(n484), .Z(n5463) );
  HS65_LL_NAND2X7 U11466 ( .A(n234), .B(n267), .Z(n5348) );
  HS65_LL_NAND2X7 U11467 ( .A(n276), .B(n309), .Z(n7055) );
  HS65_LL_NAND2X7 U11468 ( .A(n63), .B(n81), .Z(n6940) );
  HS65_LL_NAND2X7 U11469 ( .A(n503), .B(n520), .Z(n6825) );
  HS65_LL_NAND2X7 U11470 ( .A(n679), .B(n696), .Z(n5233) );
  HS65_LL_NAND2X7 U11471 ( .A(n866), .B(n848), .Z(n1352) );
  HS65_LL_NAND2X7 U11472 ( .A(n784), .B(n766), .Z(n2104) );
  HS65_LL_NAND2X7 U11473 ( .A(n825), .B(n807), .Z(n1728) );
  HS65_LL_NAND2X7 U11474 ( .A(n655), .B(n628), .Z(n3685) );
  HS65_LL_NAND2X7 U11475 ( .A(n340), .B(n325), .Z(n8586) );
  HS65_LL_NAND2X7 U11476 ( .A(n804), .B(n832), .Z(n1646) );
  HS65_LL_NAND2X7 U11477 ( .A(n438), .B(n417), .Z(n3785) );
  HS65_LL_NAND2X7 U11478 ( .A(n214), .B(n194), .Z(n3427) );
  HS65_LL_NAND4ABX3 U11479 ( .A(n8036), .B(n8500), .C(n8367), .D(n8569), .Z(
        n8889) );
  HS65_LL_NAND2X7 U11480 ( .A(n198), .B(n216), .Z(n3525) );
  HS65_LL_NAND2X7 U11481 ( .A(n886), .B(n914), .Z(n2398) );
  HS65_LL_NAND2X7 U11482 ( .A(n763), .B(n791), .Z(n2022) );
  HS65_LL_NAND2X7 U11483 ( .A(n845), .B(n873), .Z(n1270) );
  HS65_LL_NAND2X7 U11484 ( .A(n893), .B(n911), .Z(n2401) );
  HS65_LL_NAND2X7 U11485 ( .A(n811), .B(n829), .Z(n1649) );
  HS65_LL_NAND2X7 U11486 ( .A(n770), .B(n788), .Z(n2025) );
  HS65_LL_NAND2X7 U11487 ( .A(n852), .B(n870), .Z(n1273) );
  HS65_LL_NAND2X7 U11488 ( .A(n540), .B(n562), .Z(n6654) );
  HS65_LL_NAND2X7 U11489 ( .A(n18), .B(n40), .Z(n5061) );
  HS65_LL_OAI21X3 U11490 ( .A(n874), .B(n867), .C(n847), .Z(n1181) );
  HS65_LL_OAI21X3 U11491 ( .A(n792), .B(n785), .C(n765), .Z(n1933) );
  HS65_LL_NAND2X7 U11492 ( .A(n591), .B(n611), .Z(n7796) );
  HS65_LL_NAND2X7 U11493 ( .A(n111), .B(n131), .Z(n7895) );
  HS65_LL_NAND2X7 U11494 ( .A(n655), .B(n635), .Z(n3670) );
  HS65_LL_OAI21X3 U11495 ( .A(n915), .B(n908), .C(n888), .Z(n2309) );
  HS65_LL_OAI21X3 U11496 ( .A(n833), .B(n826), .C(n806), .Z(n1557) );
  HS65_LL_NAND2X7 U11497 ( .A(n497), .B(n519), .Z(n6776) );
  HS65_LL_NAND2X7 U11498 ( .A(n673), .B(n695), .Z(n5184) );
  HS65_LL_NAND2X7 U11499 ( .A(n454), .B(n482), .Z(n5415) );
  HS65_LL_NAND2X7 U11500 ( .A(n279), .B(n307), .Z(n7007) );
  HS65_LL_NAND2X7 U11501 ( .A(n237), .B(n265), .Z(n5300) );
  HS65_LL_NAND2X7 U11502 ( .A(n58), .B(n79), .Z(n6892) );
  HS65_LL_NAND2X7 U11503 ( .A(n236), .B(n265), .Z(n5277) );
  HS65_LL_NAND2X7 U11504 ( .A(n59), .B(n79), .Z(n6869) );
  HS65_LL_NAND2X7 U11505 ( .A(n761), .B(n792), .Z(n1938) );
  HS65_LL_NAND2X7 U11506 ( .A(n843), .B(n874), .Z(n1186) );
  HS65_LL_NAND2X7 U11507 ( .A(n332), .B(n347), .Z(n8547) );
  HS65_LL_NAND2X7 U11508 ( .A(n343), .B(n334), .Z(n8336) );
  HS65_LL_NAND2X7 U11509 ( .A(n884), .B(n915), .Z(n2314) );
  HS65_LL_NAND2X7 U11510 ( .A(n261), .B(n235), .Z(n5347) );
  HS65_LL_NAND2X7 U11511 ( .A(n303), .B(n277), .Z(n7054) );
  HS65_LL_NAND2X7 U11512 ( .A(n85), .B(n66), .Z(n6939) );
  HS65_LL_NAND2X7 U11513 ( .A(n802), .B(n833), .Z(n1562) );
  HS65_LL_NAND4ABX3 U11514 ( .A(n1962), .B(n1963), .C(n1964), .D(n1965), .Z(
        n1923) );
  HS65_LL_NAND4ABX3 U11515 ( .A(n1991), .B(n1992), .C(n1993), .D(n1994), .Z(
        n1963) );
  HS65_LL_NOR4ABX2 U11516 ( .A(n1966), .B(n1967), .C(n1968), .D(n1969), .Z(
        n1965) );
  HS65_LL_MX41X7 U11517 ( .D0(n782), .S0(n763), .D1(n793), .S1(n760), .D2(n778), .S2(n768), .D3(n790), .S3(n765), .Z(n1962) );
  HS65_LL_NAND4ABX3 U11518 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .Z(
        n1171) );
  HS65_LL_NAND4ABX3 U11519 ( .A(n1239), .B(n1240), .C(n1241), .D(n1242), .Z(
        n1211) );
  HS65_LL_NOR4ABX2 U11520 ( .A(n1214), .B(n1215), .C(n1216), .D(n1217), .Z(
        n1213) );
  HS65_LL_MX41X7 U11521 ( .D0(n864), .S0(n845), .D1(n875), .S1(n842), .D2(n860), .S2(n850), .D3(n872), .S3(n847), .Z(n1210) );
  HS65_LL_NAND2X7 U11522 ( .A(n431), .B(n406), .Z(n3176) );
  HS65_LL_NAND2X7 U11523 ( .A(n225), .B(n203), .Z(n2949) );
  HS65_LL_NAND4ABX3 U11524 ( .A(n2338), .B(n2339), .C(n2340), .D(n2341), .Z(
        n2299) );
  HS65_LL_NAND4ABX3 U11525 ( .A(n2367), .B(n2368), .C(n2369), .D(n2370), .Z(
        n2339) );
  HS65_LL_MX41X7 U11526 ( .D0(n905), .S0(n886), .D1(n916), .S1(n883), .D2(n901), .S2(n891), .D3(n913), .S3(n888), .Z(n2338) );
  HS65_LL_NOR4ABX2 U11527 ( .A(n2342), .B(n2343), .C(n2344), .D(n2345), .Z(
        n2341) );
  HS65_LL_NAND4ABX3 U11528 ( .A(n1586), .B(n1587), .C(n1588), .D(n1589), .Z(
        n1547) );
  HS65_LL_NOR4ABX2 U11529 ( .A(n1590), .B(n1591), .C(n1592), .D(n1593), .Z(
        n1589) );
  HS65_LL_NAND4ABX3 U11530 ( .A(n1615), .B(n1616), .C(n1617), .D(n1618), .Z(
        n1587) );
  HS65_LL_MX41X7 U11531 ( .D0(n823), .S0(n804), .D1(n834), .S1(n801), .D2(n819), .S2(n809), .D3(n831), .S3(n806), .Z(n1586) );
  HS65_LL_NAND2X7 U11532 ( .A(n885), .B(n902), .Z(n2446) );
  HS65_LL_NAND2X7 U11533 ( .A(n762), .B(n779), .Z(n2070) );
  HS65_LL_NAND2X7 U11534 ( .A(n413), .B(n436), .Z(n3879) );
  HS65_LL_NAND2X7 U11535 ( .A(n644), .B(n625), .Z(n3150) );
  HS65_LL_NAND2X7 U11536 ( .A(n353), .B(n328), .Z(n8331) );
  HS65_LL_NAND2X7 U11537 ( .A(n247), .B(n265), .Z(n4919) );
  HS65_LL_NAND2X7 U11538 ( .A(n68), .B(n79), .Z(n6512) );
  HS65_LL_NAND2X7 U11539 ( .A(n289), .B(n307), .Z(n6565) );
  HS65_LL_NAND2X7 U11540 ( .A(n844), .B(n861), .Z(n1318) );
  HS65_LL_NAND2X7 U11541 ( .A(n803), .B(n820), .Z(n1694) );
  HS65_LL_IVX9 U11542 ( .A(n2796), .Z(n231) );
  HS65_LL_IVX9 U11543 ( .A(n2788), .Z(n53) );
  HS65_LL_OAI21X3 U11544 ( .A(n369), .B(n362), .C(n396), .Z(n8650) );
  HS65_LL_NAND2X7 U11545 ( .A(n823), .B(n800), .Z(n1566) );
  HS65_LL_NAND2X7 U11546 ( .A(n864), .B(n841), .Z(n1190) );
  HS65_LL_NAND2X7 U11547 ( .A(n782), .B(n759), .Z(n1942) );
  HS65_LL_NAND2X7 U11548 ( .A(n650), .B(n628), .Z(n3730) );
  HS65_LLS_XOR3X2 U11549 ( .A(n2659), .B(n2654), .C(n2660), .Z(n2658) );
  HS65_LL_NAND2X7 U11550 ( .A(n905), .B(n882), .Z(n2318) );
  HS65_LL_NAND2X7 U11551 ( .A(n441), .B(n409), .Z(n3845) );
  HS65_LL_NAND2X7 U11552 ( .A(n888), .B(n905), .Z(n2457) );
  HS65_LL_NAND2X7 U11553 ( .A(n765), .B(n782), .Z(n2081) );
  HS65_LL_NAND2X7 U11554 ( .A(n847), .B(n864), .Z(n1329) );
  HS65_LL_NAND2X7 U11555 ( .A(n806), .B(n823), .Z(n1705) );
  HS65_LL_NAND2X7 U11556 ( .A(n658), .B(n637), .Z(n3741) );
  HS65_LL_NAND2X7 U11557 ( .A(n427), .B(n419), .Z(n3856) );
  HS65_LL_NAND2X7 U11558 ( .A(n614), .B(n590), .Z(n8711) );
  HS65_LL_NAND2X7 U11559 ( .A(n134), .B(n110), .Z(n8801) );
  HS65_LL_NAND2X7 U11560 ( .A(n766), .B(n779), .Z(n2122) );
  HS65_LL_NAND2X7 U11561 ( .A(n848), .B(n861), .Z(n1370) );
  HS65_LL_NAND2X7 U11562 ( .A(n785), .B(n771), .Z(n2061) );
  HS65_LL_NAND2X7 U11563 ( .A(n867), .B(n853), .Z(n1309) );
  HS65_LL_NAND2X7 U11564 ( .A(n209), .B(n191), .Z(n3501) );
  HS65_LL_NAND2X7 U11565 ( .A(n889), .B(n902), .Z(n2498) );
  HS65_LL_NAND2X7 U11566 ( .A(n826), .B(n812), .Z(n1685) );
  HS65_LL_NAND2X7 U11567 ( .A(n908), .B(n894), .Z(n2437) );
  HS65_LL_NAND2X7 U11568 ( .A(n807), .B(n820), .Z(n1746) );
  HS65_LL_NAND2X7 U11569 ( .A(n564), .B(n536), .Z(n6675) );
  HS65_LL_NAND2X7 U11570 ( .A(n42), .B(n14), .Z(n5082) );
  HS65_LL_NAND2X7 U11571 ( .A(n395), .B(n365), .Z(n8099) );
  HS65_LL_NAND2X7 U11572 ( .A(n395), .B(n376), .Z(n8098) );
  HS65_LL_NAND2X7 U11573 ( .A(n353), .B(n319), .Z(n8332) );
  HS65_LL_NAND2X7 U11574 ( .A(n374), .B(n383), .Z(n8245) );
  HS65_LL_NAND2X7 U11575 ( .A(n341), .B(n329), .Z(n8587) );
  HS65_LL_NAND2X7 U11576 ( .A(n267), .B(n240), .Z(n5304) );
  HS65_LL_NAND2X7 U11577 ( .A(n484), .B(n457), .Z(n5419) );
  HS65_LL_NAND2X7 U11578 ( .A(n696), .B(n676), .Z(n5188) );
  HS65_LL_NAND2X7 U11579 ( .A(n81), .B(n62), .Z(n6896) );
  HS65_LL_NAND2X7 U11580 ( .A(n309), .B(n282), .Z(n7011) );
  HS65_LL_NAND2X7 U11581 ( .A(n520), .B(n500), .Z(n6780) );
  HS65_LL_NAND2X7 U11582 ( .A(n41), .B(n21), .Z(n5066) );
  HS65_LL_NAND2X7 U11583 ( .A(n563), .B(n543), .Z(n6659) );
  HS65_LL_NAND2X7 U11584 ( .A(n391), .B(n377), .Z(n8285) );
  HS65_LLS_XOR3X2 U11585 ( .A(n7546), .B(n2618), .C(n2751), .Z(n7559) );
  HS65_LL_NAND2X7 U11586 ( .A(n864), .B(n844), .Z(n1230) );
  HS65_LL_NAND2X7 U11587 ( .A(n782), .B(n762), .Z(n1982) );
  HS65_LL_NAND2X7 U11588 ( .A(n905), .B(n885), .Z(n2358) );
  HS65_LL_NAND2X7 U11589 ( .A(n823), .B(n803), .Z(n1606) );
  HS65_LL_NAND2X7 U11590 ( .A(n41), .B(n24), .Z(n5097) );
  HS65_LL_NAND2X7 U11591 ( .A(n563), .B(n546), .Z(n6690) );
  HS65_LL_NAND2X7 U11592 ( .A(n660), .B(n628), .Z(n3764) );
  HS65_LL_OAI21X3 U11593 ( .A(n825), .B(n1594), .C(n799), .Z(n1591) );
  HS65_LL_NAND2X7 U11594 ( .A(n599), .B(n578), .Z(n8682) );
  HS65_LL_NAND2X7 U11595 ( .A(n119), .B(n98), .Z(n8772) );
  HS65_LL_OAI21X3 U11596 ( .A(n907), .B(n2346), .C(n881), .Z(n2343) );
  HS65_LL_OAI21X3 U11597 ( .A(n784), .B(n1970), .C(n758), .Z(n1967) );
  HS65_LL_OAI21X3 U11598 ( .A(n866), .B(n1218), .C(n840), .Z(n1215) );
  HS65_LL_NAND2X7 U11599 ( .A(n324), .B(n344), .Z(n8588) );
  HS65_LL_NAND2X7 U11600 ( .A(n531), .B(n559), .Z(n6673) );
  HS65_LL_NAND2X7 U11601 ( .A(n9), .B(n37), .Z(n5080) );
  HS65_LL_NOR4ABX2 U11602 ( .A(n1843), .B(n1728), .C(n1616), .D(n1647), .Z(
        n1837) );
  HS65_LL_OAI21X3 U11603 ( .A(n822), .B(n823), .C(n813), .Z(n1843) );
  HS65_LL_NAND2X7 U11604 ( .A(n699), .B(n670), .Z(n5144) );
  HS65_LL_NAND2X7 U11605 ( .A(n523), .B(n494), .Z(n6736) );
  HS65_LL_NAND2X7 U11606 ( .A(n90), .B(n55), .Z(n6853) );
  HS65_LL_NAND2X7 U11607 ( .A(n255), .B(n244), .Z(n5261) );
  HS65_LL_NAND2X7 U11608 ( .A(n472), .B(n461), .Z(n5376) );
  HS65_LL_NAND2X7 U11609 ( .A(n297), .B(n286), .Z(n6968) );
  HS65_LL_NAND2X7 U11610 ( .A(n333), .B(n349), .Z(n8359) );
  HS65_LL_NAND2X7 U11611 ( .A(n320), .B(n342), .Z(n8551) );
  HS65_LL_NAND2X7 U11612 ( .A(n82), .B(n68), .Z(n6849) );
  HS65_LL_NAND2X7 U11613 ( .A(n268), .B(n247), .Z(n5257) );
  HS65_LL_NAND2X7 U11614 ( .A(n485), .B(n464), .Z(n5372) );
  HS65_LL_NAND2X7 U11615 ( .A(n310), .B(n289), .Z(n6964) );
  HS65_LL_NAND2X7 U11616 ( .A(n518), .B(n490), .Z(n6732) );
  HS65_LL_NAND2X7 U11617 ( .A(n124), .B(n100), .Z(n7922) );
  HS65_LL_NAND2X7 U11618 ( .A(n604), .B(n580), .Z(n7824) );
  HS65_LL_NAND4ABX3 U11619 ( .A(n6121), .B(n6122), .C(n6123), .D(n6124), .Z(
        n6111) );
  HS65_LL_AOI212X4 U11620 ( .A(n494), .B(n512), .C(n490), .D(n526), .E(n6125), 
        .Z(n6124) );
  HS65_LL_NAND4ABX3 U11621 ( .A(n4528), .B(n4529), .C(n4530), .D(n4531), .Z(
        n4518) );
  HS65_LL_AOI212X4 U11622 ( .A(n670), .B(n688), .C(n666), .D(n702), .E(n4532), 
        .Z(n4531) );
  HS65_LL_NOR2X6 U11623 ( .A(n788), .B(n785), .Z(n2118) );
  HS65_LL_NOR2X6 U11624 ( .A(n870), .B(n867), .Z(n1366) );
  HS65_LL_NOR2X6 U11625 ( .A(n911), .B(n908), .Z(n2494) );
  HS65_LL_NOR2X6 U11626 ( .A(n829), .B(n826), .Z(n1742) );
  HS65_LL_NAND2X7 U11627 ( .A(n367), .B(n394), .Z(n8253) );
  HS65_LLS_XNOR2X6 U11628 ( .A(n2687), .B(n2627), .Z(n2636) );
  HS65_LL_NAND2X7 U11629 ( .A(n627), .B(n645), .Z(n3723) );
  HS65_LL_NAND2X7 U11630 ( .A(n890), .B(n902), .Z(n2484) );
  HS65_LL_NAND2X7 U11631 ( .A(n849), .B(n861), .Z(n1356) );
  HS65_LL_NAND2X7 U11632 ( .A(n767), .B(n779), .Z(n2108) );
  HS65_LL_NAND2X7 U11633 ( .A(n369), .B(n383), .Z(n8267) );
  HS65_LL_NAND2X7 U11634 ( .A(n808), .B(n820), .Z(n1732) );
  HS65_LL_NAND2X7 U11635 ( .A(n440), .B(n409), .Z(n3883) );
  HS65_LL_AOI12X2 U11636 ( .A(n156), .B(n164), .C(n3651), .Z(n3648) );
  HS65_LL_NOR2X6 U11637 ( .A(n869), .B(n1260), .Z(n1316) );
  HS65_LL_NOR2X6 U11638 ( .A(n787), .B(n2012), .Z(n2068) );
  HS65_LL_NOR2X6 U11639 ( .A(n910), .B(n2388), .Z(n2444) );
  HS65_LL_NOR2X6 U11640 ( .A(n828), .B(n1636), .Z(n1692) );
  HS65_LL_NOR2X6 U11641 ( .A(n416), .B(n3775), .Z(n3844) );
  HS65_LL_NOR2X6 U11642 ( .A(n54), .B(n6832), .Z(n6856) );
  HS65_LL_NOR2X6 U11643 ( .A(n242), .B(n5240), .Z(n5264) );
  HS65_LL_AOI12X2 U11644 ( .A(n907), .B(n891), .C(n2462), .Z(n2459) );
  HS65_LL_AOI12X2 U11645 ( .A(n784), .B(n768), .C(n2086), .Z(n2083) );
  HS65_LL_AOI12X2 U11646 ( .A(n866), .B(n850), .C(n1334), .Z(n1331) );
  HS65_LL_AOI12X2 U11647 ( .A(n825), .B(n809), .C(n1710), .Z(n1707) );
  HS65_LL_AOI12X2 U11648 ( .A(n413), .B(n435), .C(n3861), .Z(n3858) );
  HS65_LL_AOI12X2 U11649 ( .A(n198), .B(n223), .C(n3507), .Z(n3504) );
  HS65_LL_AOI12X2 U11650 ( .A(n631), .B(n648), .C(n3746), .Z(n3743) );
  HS65_LL_NAND2X7 U11651 ( .A(n367), .B(n398), .Z(n8074) );
  HS65_LL_AOI12X2 U11652 ( .A(n167), .B(n151), .C(n3543), .Z(n4149) );
  HS65_LL_NAND4ABX3 U11653 ( .A(n1276), .B(n1372), .C(n1443), .D(n1251), .Z(
        n1439) );
  HS65_LL_OAI21X3 U11654 ( .A(n873), .B(n865), .C(n850), .Z(n1443) );
  HS65_LL_NAND4ABX3 U11655 ( .A(n2028), .B(n2124), .C(n2195), .D(n2003), .Z(
        n2191) );
  HS65_LL_OAI21X3 U11656 ( .A(n791), .B(n783), .C(n768), .Z(n2195) );
  HS65_LL_NAND4ABX3 U11657 ( .A(n1652), .B(n1748), .C(n1819), .D(n1627), .Z(
        n1815) );
  HS65_LL_OAI21X3 U11658 ( .A(n832), .B(n824), .C(n809), .Z(n1819) );
  HS65_LL_AO212X4 U11659 ( .A(n869), .B(n1300), .C(n870), .D(n851), .E(n1473), 
        .Z(n1472) );
  HS65_LL_CB4I6X9 U11660 ( .A(n871), .B(n872), .C(n850), .D(n1373), .Z(n1473)
         );
  HS65_LL_AO212X4 U11661 ( .A(n787), .B(n2052), .C(n788), .D(n769), .E(n2225), 
        .Z(n2224) );
  HS65_LL_CB4I6X9 U11662 ( .A(n789), .B(n790), .C(n768), .D(n2125), .Z(n2225)
         );
  HS65_LL_AO212X4 U11663 ( .A(n828), .B(n1676), .C(n829), .D(n810), .E(n1849), 
        .Z(n1848) );
  HS65_LL_CB4I6X9 U11664 ( .A(n830), .B(n831), .C(n809), .D(n1749), .Z(n1849)
         );
  HS65_LL_AO212X4 U11665 ( .A(n910), .B(n2428), .C(n911), .D(n892), .E(n2601), 
        .Z(n2600) );
  HS65_LL_CB4I6X9 U11666 ( .A(n912), .B(n913), .C(n891), .D(n2501), .Z(n2601)
         );
  HS65_LL_AO212X4 U11667 ( .A(n416), .B(n434), .C(n412), .D(n428), .E(n4336), 
        .Z(n4335) );
  HS65_LL_CB4I6X9 U11668 ( .A(n407), .B(n411), .C(n435), .D(n3802), .Z(n4336)
         );
  HS65_LL_NAND4ABX3 U11669 ( .A(n6860), .B(n6861), .C(n6862), .D(n6863), .Z(
        n6845) );
  HS65_LL_NAND4ABX3 U11670 ( .A(n5268), .B(n5269), .C(n5270), .D(n5271), .Z(
        n5253) );
  HS65_LL_NAND4ABX3 U11671 ( .A(n2040), .B(n2041), .C(n2042), .D(n2043), .Z(
        n2034) );
  HS65_LL_NAND4ABX3 U11672 ( .A(n1288), .B(n1289), .C(n1290), .D(n1291), .Z(
        n1282) );
  HS65_LL_NAND4ABX3 U11673 ( .A(n1664), .B(n1665), .C(n1666), .D(n1667), .Z(
        n1658) );
  HS65_LL_NAND4ABX3 U11674 ( .A(n2416), .B(n2417), .C(n2418), .D(n2419), .Z(
        n2410) );
  HS65_LL_NAND4ABX3 U11675 ( .A(n3747), .B(n3748), .C(n3749), .D(n3750), .Z(
        n3737) );
  HS65_LL_NAND4ABX3 U11676 ( .A(n1715), .B(n1716), .C(n1717), .D(n1718), .Z(
        n1700) );
  HS65_LL_NAND4ABX3 U11677 ( .A(n1339), .B(n1340), .C(n1341), .D(n1342), .Z(
        n1324) );
  HS65_LL_NAND4ABX3 U11678 ( .A(n2091), .B(n2092), .C(n2093), .D(n2094), .Z(
        n2076) );
  HS65_LL_NAND4ABX3 U11679 ( .A(n2467), .B(n2468), .C(n2469), .D(n2470), .Z(
        n2452) );
  HS65_LL_NAND4ABX3 U11680 ( .A(n3512), .B(n3513), .C(n3514), .D(n3515), .Z(
        n3496) );
  HS65_LL_NAND3AX6 U11681 ( .A(n1986), .B(n1987), .C(n1988), .Z(n1973) );
  HS65_LL_AOI12X2 U11682 ( .A(n786), .B(n1989), .C(n1990), .Z(n1988) );
  HS65_LL_NAND3AX6 U11683 ( .A(n1234), .B(n1235), .C(n1236), .Z(n1221) );
  HS65_LL_AOI12X2 U11684 ( .A(n868), .B(n1237), .C(n1238), .Z(n1236) );
  HS65_LL_NAND4ABX3 U11685 ( .A(n4946), .B(n5445), .C(n4985), .D(n5912), .Z(
        n5906) );
  HS65_LL_OAI21X3 U11686 ( .A(n484), .B(n479), .C(n464), .Z(n5912) );
  HS65_LL_NAND4ABX3 U11687 ( .A(n6539), .B(n7037), .C(n6578), .D(n7504), .Z(
        n7498) );
  HS65_LL_OAI21X3 U11688 ( .A(n309), .B(n304), .C(n289), .Z(n7504) );
  HS65_LL_NAND4ABX3 U11689 ( .A(n4893), .B(n5330), .C(n4932), .D(n5853), .Z(
        n5847) );
  HS65_LL_OAI21X3 U11690 ( .A(n267), .B(n262), .C(n247), .Z(n5853) );
  HS65_LL_NAND4ABX3 U11691 ( .A(n6486), .B(n6922), .C(n6525), .D(n7445), .Z(
        n7439) );
  HS65_LL_OAI21X3 U11692 ( .A(n81), .B(n84), .C(n68), .Z(n7445) );
  HS65_LL_NAND3AX6 U11693 ( .A(n2362), .B(n2363), .C(n2364), .Z(n2349) );
  HS65_LL_AOI12X2 U11694 ( .A(n909), .B(n2365), .C(n2366), .Z(n2364) );
  HS65_LL_NAND4ABX3 U11695 ( .A(n8409), .B(n8401), .C(n8740), .D(n9026), .Z(
        n9022) );
  HS65_LL_OAI21X3 U11696 ( .A(n610), .B(n606), .C(n583), .Z(n9026) );
  HS65_LL_NAND4ABX3 U11697 ( .A(n8461), .B(n8453), .C(n8830), .D(n9084), .Z(
        n9080) );
  HS65_LL_OAI21X3 U11698 ( .A(n130), .B(n126), .C(n103), .Z(n9084) );
  HS65_LL_IVX9 U11699 ( .A(n2758), .Z(n529) );
  HS65_LL_NAND3AX6 U11700 ( .A(n8270), .B(n8271), .C(n8272), .Z(n8259) );
  HS65_LL_AOI12X2 U11701 ( .A(n378), .B(n386), .C(n8273), .Z(n8272) );
  HS65_LL_NAND4ABX3 U11702 ( .A(n3862), .B(n3863), .C(n3864), .D(n3865), .Z(
        n3852) );
  HS65_LL_NAND3X5 U11703 ( .A(n1653), .B(n1654), .C(n1655), .Z(n1641) );
  HS65_LL_AOI12X2 U11704 ( .A(n811), .B(n828), .C(n1656), .Z(n1655) );
  HS65_LL_IVX9 U11705 ( .A(n2782), .Z(n50) );
  HS65_LL_NAND4ABX3 U11706 ( .A(n2448), .B(n2449), .C(n2450), .D(n2451), .Z(
        n2433) );
  HS65_LL_NAND4ABX3 U11707 ( .A(n1320), .B(n1321), .C(n1322), .D(n1323), .Z(
        n1305) );
  HS65_LL_NAND4ABX3 U11708 ( .A(n2072), .B(n2073), .C(n2074), .D(n2075), .Z(
        n2057) );
  HS65_LL_NAND4ABX3 U11709 ( .A(n4991), .B(n5397), .C(n4798), .D(n5358), .Z(
        n5918) );
  HS65_LL_NAND4ABX3 U11710 ( .A(n6584), .B(n6989), .C(n6391), .D(n6950), .Z(
        n7510) );
  HS65_LL_NAND4ABX3 U11711 ( .A(n4879), .B(n5282), .C(n4737), .D(n5243), .Z(
        n5859) );
  HS65_LL_NAND4ABX3 U11712 ( .A(n6472), .B(n6874), .C(n6352), .D(n6835), .Z(
        n7451) );
  HS65_LL_NAND4ABX3 U11713 ( .A(n4865), .B(n5165), .C(n4652), .D(n5125), .Z(
        n5787) );
  HS65_LL_NAND4ABX3 U11714 ( .A(n6458), .B(n6757), .C(n6245), .D(n6717), .Z(
        n7379) );
  HS65_LL_NAND4ABX3 U11715 ( .A(n8418), .B(n8133), .C(n8669), .D(n8697), .Z(
        n9008) );
  HS65_LL_NAND4ABX3 U11716 ( .A(n8470), .B(n8184), .C(n8759), .D(n8787), .Z(
        n9066) );
  HS65_LL_MX41X7 U11717 ( .D0(n864), .S0(n848), .D1(n868), .S1(n849), .D2(n865), .S2(n843), .D3(n860), .S3(n844), .Z(n1422) );
  HS65_LL_NAND4ABX3 U11718 ( .A(n6595), .B(n6166), .C(n6258), .D(n6635), .Z(
        n7317) );
  HS65_LL_NAND4ABX3 U11719 ( .A(n5002), .B(n4573), .C(n4665), .D(n5042), .Z(
        n5725) );
  HS65_LL_MX41X7 U11720 ( .D0(n165), .S0(n143), .D1(n153), .S1(n164), .D2(n154), .S2(n172), .D3(n163), .S3(n151), .Z(n4129) );
  HS65_LL_MX41X7 U11721 ( .D0(n793), .S0(n767), .D1(n784), .S1(n772), .D2(n765), .S2(n788), .D3(n758), .S3(n779), .Z(n2162) );
  HS65_LL_MX41X7 U11722 ( .D0(n865), .S0(n843), .D1(n867), .S1(n850), .D2(n860), .S2(n853), .D3(n844), .S3(n874), .Z(n1256) );
  HS65_LL_MX41X7 U11723 ( .D0(n875), .S0(n849), .D1(n866), .S1(n854), .D2(n847), .S2(n870), .D3(n840), .S3(n861), .Z(n1410) );
  HS65_LL_MX41X7 U11724 ( .D0(n834), .S0(n808), .D1(n825), .S1(n813), .D2(n806), .S2(n829), .D3(n799), .S3(n820), .Z(n1786) );
  HS65_LL_MX41X7 U11725 ( .D0(n916), .S0(n890), .D1(n907), .S1(n895), .D2(n888), .S2(n911), .D3(n881), .S3(n902), .Z(n2538) );
  HS65_LL_MX41X7 U11726 ( .D0(n916), .S0(n881), .D1(n883), .S1(n911), .D2(n892), .S2(n902), .D3(n913), .S3(n882), .Z(n2578) );
  HS65_LL_MX41X7 U11727 ( .D0(n793), .S0(n758), .D1(n760), .S1(n788), .D2(n769), .S2(n779), .D3(n790), .S3(n759), .Z(n2202) );
  HS65_LL_MX41X7 U11728 ( .D0(n875), .S0(n840), .D1(n842), .S1(n870), .D2(n851), .S2(n861), .D3(n872), .S3(n841), .Z(n1450) );
  HS65_LL_MX41X7 U11729 ( .D0(n834), .S0(n799), .D1(n801), .S1(n829), .D2(n810), .S2(n820), .D3(n831), .S3(n800), .Z(n1826) );
  HS65_LL_MX41X7 U11730 ( .D0(n781), .S0(n769), .D1(n778), .S1(n757), .D2(n758), .S2(n791), .D3(n759), .S3(n789), .Z(n2018) );
  HS65_LL_MX41X7 U11731 ( .D0(n904), .S0(n892), .D1(n901), .S1(n880), .D2(n881), .S2(n914), .D3(n882), .S3(n912), .Z(n2394) );
  HS65_LL_MX41X7 U11732 ( .D0(n863), .S0(n851), .D1(n860), .S1(n839), .D2(n840), .S2(n873), .D3(n841), .S3(n871), .Z(n1266) );
  HS65_LL_MX41X7 U11733 ( .D0(n418), .S0(n428), .D1(n405), .S1(n433), .D2(n443), .S2(n417), .D3(n439), .S3(n407), .Z(n3781) );
  HS65_LL_MX41X7 U11734 ( .D0(n636), .S0(n659), .D1(n624), .S1(n646), .D2(n652), .S2(n635), .D3(n656), .S3(n626), .Z(n3666) );
  HS65_LL_AND3X9 U11735 ( .A(n2196), .B(n2197), .C(n2198), .Z(n2140) );
  HS65_LL_NOR4X4 U11736 ( .A(n1980), .B(n1991), .C(n1999), .D(n2040), .Z(n2197) );
  HS65_LL_NOR4ABX2 U11737 ( .A(n2051), .B(n1902), .C(n2063), .D(n2115), .Z(
        n2196) );
  HS65_LL_NOR4ABX2 U11738 ( .A(n2199), .B(n1938), .C(n2106), .D(n2200), .Z(
        n2198) );
  HS65_LL_AND3X9 U11739 ( .A(n1444), .B(n1445), .C(n1446), .Z(n1388) );
  HS65_LL_NOR4X4 U11740 ( .A(n1228), .B(n1239), .C(n1247), .D(n1288), .Z(n1445) );
  HS65_LL_NOR4ABX2 U11741 ( .A(n1299), .B(n1150), .C(n1311), .D(n1363), .Z(
        n1444) );
  HS65_LL_NOR4ABX2 U11742 ( .A(n1447), .B(n1186), .C(n1354), .D(n1448), .Z(
        n1446) );
  HS65_LL_AND3X9 U11743 ( .A(n1820), .B(n1821), .C(n1822), .Z(n1764) );
  HS65_LL_NOR4X4 U11744 ( .A(n1604), .B(n1615), .C(n1623), .D(n1664), .Z(n1821) );
  HS65_LL_NOR4ABX2 U11745 ( .A(n1675), .B(n1526), .C(n1687), .D(n1739), .Z(
        n1820) );
  HS65_LL_NOR4ABX2 U11746 ( .A(n1823), .B(n1562), .C(n1730), .D(n1824), .Z(
        n1822) );
  HS65_LL_AND3X9 U11747 ( .A(n2572), .B(n2573), .C(n2574), .Z(n2516) );
  HS65_LL_NOR4X4 U11748 ( .A(n2356), .B(n2367), .C(n2375), .D(n2416), .Z(n2573) );
  HS65_LL_NOR4ABX2 U11749 ( .A(n2427), .B(n2278), .C(n2439), .D(n2491), .Z(
        n2572) );
  HS65_LL_NOR4ABX2 U11750 ( .A(n2575), .B(n2314), .C(n2482), .D(n2576), .Z(
        n2574) );
  HS65_LL_AND3X9 U11751 ( .A(n4204), .B(n4205), .C(n4206), .Z(n4064) );
  HS65_LL_NOR4X4 U11752 ( .A(n3090), .B(n3103), .C(n3117), .D(n3457), .Z(n4205) );
  HS65_LL_NOR4ABX2 U11753 ( .A(n3472), .B(n2862), .C(n3484), .D(n3445), .Z(
        n4204) );
  HS65_LL_NOR4ABX2 U11754 ( .A(n4207), .B(n2949), .C(n3527), .D(n4208), .Z(
        n4206) );
  HS65_LL_AND3X9 U11755 ( .A(n4307), .B(n4308), .C(n4309), .Z(n3966) );
  HS65_LL_NOR4X4 U11756 ( .A(n3375), .B(n3386), .C(n3398), .D(n3814), .Z(n4308) );
  HS65_LL_NOR4ABX2 U11757 ( .A(n3828), .B(n2999), .C(n3839), .D(n3803), .Z(
        n4307) );
  HS65_LL_NOR4ABX2 U11758 ( .A(n4310), .B(n3176), .C(n3881), .D(n4311), .Z(
        n4309) );
  HS65_LL_AND3X9 U11759 ( .A(n4248), .B(n4249), .C(n4250), .Z(n3946) );
  HS65_LL_NOR4X4 U11760 ( .A(n3321), .B(n3332), .C(n3344), .D(n3699), .Z(n4249) );
  HS65_LL_NOR4ABX2 U11761 ( .A(n3764), .B(n3150), .C(n4251), .D(n4252), .Z(
        n4250) );
  HS65_LL_NOR4ABX2 U11762 ( .A(n3713), .B(n2974), .C(n3725), .D(n3688), .Z(
        n4248) );
  HS65_LL_CBI4I6X5 U11763 ( .A(n847), .B(n1300), .C(n867), .D(n1395), .Z(n1375) );
  HS65_LL_OA12X9 U11764 ( .A(n1218), .B(n872), .C(n851), .Z(n1395) );
  HS65_LL_OA12X9 U11765 ( .A(n1989), .B(n770), .C(n793), .Z(n2161) );
  HS65_LL_OA12X9 U11766 ( .A(n1237), .B(n852), .C(n875), .Z(n1409) );
  HS65_LL_OA12X9 U11767 ( .A(n1613), .B(n811), .C(n834), .Z(n1785) );
  HS65_LL_OA12X9 U11768 ( .A(n2365), .B(n893), .C(n916), .Z(n2537) );
  HS65_LL_NAND3X5 U11769 ( .A(n9005), .B(n9006), .C(n9007), .Z(n7698) );
  HS65_LL_NOR4ABX2 U11770 ( .A(n8682), .B(n8003), .C(n8716), .D(n8738), .Z(
        n9005) );
  HS65_LL_NOR4ABX2 U11771 ( .A(n8403), .B(n8408), .C(n8749), .D(n8393), .Z(
        n9006) );
  HS65_LL_NOR4X4 U11772 ( .A(n8712), .B(n8152), .C(n9008), .D(n9009), .Z(n9007) );
  HS65_LL_NAND3X5 U11773 ( .A(n9063), .B(n9064), .C(n9065), .Z(n7736) );
  HS65_LL_NOR4ABX2 U11774 ( .A(n8772), .B(n8016), .C(n8806), .D(n8828), .Z(
        n9063) );
  HS65_LL_NOR4ABX2 U11775 ( .A(n8455), .B(n8460), .C(n8839), .D(n8445), .Z(
        n9064) );
  HS65_LL_NOR4X4 U11776 ( .A(n8802), .B(n8175), .C(n9066), .D(n9067), .Z(n9065) );
  HS65_LL_IVX9 U11777 ( .A(n8807), .Z(n109) );
  HS65_LL_AND3X9 U11778 ( .A(n5373), .B(n4780), .C(n5391), .Z(n5904) );
  HS65_LL_AND3X9 U11779 ( .A(n6965), .B(n6373), .C(n6983), .Z(n7496) );
  HS65_LL_AND3X9 U11780 ( .A(n5258), .B(n4753), .C(n5276), .Z(n5845) );
  HS65_LL_AND3X9 U11781 ( .A(n6850), .B(n6334), .C(n6868), .Z(n7437) );
  HS65_LLS_XNOR2X6 U11782 ( .A(n2821), .B(n2797), .Z(n4393) );
  HS65_LLS_XNOR2X6 U11783 ( .A(n2813), .B(n2789), .Z(n5986) );
  HS65_LLS_XNOR2X6 U11784 ( .A(n3213), .B(n2770), .Z(n4395) );
  HS65_LLS_XNOR2X6 U11785 ( .A(n3205), .B(n2762), .Z(n5988) );
  HS65_LLS_XNOR2X6 U11786 ( .A(n3211), .B(n2768), .Z(n4402) );
  HS65_LLS_XNOR2X6 U11787 ( .A(n3008), .B(n2760), .Z(n5995) );
  HS65_LLS_XNOR2X6 U11788 ( .A(n3003), .B(n361), .Z(n7572) );
  HS65_LLS_XNOR2X6 U11789 ( .A(n3000), .B(n2752), .Z(n7585) );
  HS65_LLS_XOR2X6 U11790 ( .A(n3533), .B(n2773), .Z(n4803) );
  HS65_LLS_XOR2X6 U11791 ( .A(n3208), .B(n2765), .Z(n6396) );
  HS65_LL_NAND4ABX3 U11792 ( .A(n6710), .B(n6711), .C(n6712), .D(n6713), .Z(
        n3009) );
  HS65_LL_MX41X7 U11793 ( .D0(n503), .S0(n521), .D1(n509), .S1(n504), .D2(n508), .S2(n501), .D3(n502), .S3(n6231), .Z(n6711) );
  HS65_LL_AOI212X4 U11794 ( .A(n519), .B(n6714), .C(n497), .D(n6447), .E(n6715), .Z(n6713) );
  HS65_LL_MX41X7 U11795 ( .D0(n493), .S0(n525), .D1(n523), .S1(n500), .D2(n526), .S2(n498), .D3(n499), .S3(n512), .Z(n6710) );
  HS65_LL_NAND4ABX3 U11796 ( .A(n6589), .B(n6590), .C(n6591), .D(n6592), .Z(
        n2761) );
  HS65_LL_MX41X7 U11797 ( .D0(n546), .S0(n564), .D1(n552), .S1(n547), .D2(n551), .S2(n544), .D3(n545), .S3(n6154), .Z(n6590) );
  HS65_LL_AOI212X4 U11798 ( .A(n562), .B(n6593), .C(n540), .D(n6309), .E(n6594), .Z(n6592) );
  HS65_LL_MX41X7 U11799 ( .D0(n536), .S0(n568), .D1(n566), .S1(n543), .D2(n569), .S2(n541), .D3(n542), .S3(n555), .Z(n6589) );
  HS65_LLS_XOR2X6 U11800 ( .A(n2802), .B(n2778), .Z(n7544) );
  HS65_LL_NAND4ABX3 U11801 ( .A(n4996), .B(n4997), .C(n4998), .D(n4999), .Z(
        n2769) );
  HS65_LL_MX41X7 U11802 ( .D0(n24), .S0(n42), .D1(n30), .S1(n25), .D2(n29), 
        .S2(n22), .D3(n23), .S3(n4561), .Z(n4997) );
  HS65_LL_AOI212X4 U11803 ( .A(n40), .B(n5000), .C(n18), .D(n4716), .E(n5001), 
        .Z(n4999) );
  HS65_LL_MX41X7 U11804 ( .D0(n14), .S0(n46), .D1(n44), .S1(n21), .D2(n47), 
        .S2(n19), .D3(n20), .S3(n33), .Z(n4996) );
  HS65_LLS_XOR2X6 U11805 ( .A(n2771), .B(n3214), .Z(n4389) );
  HS65_LLS_XOR2X6 U11806 ( .A(n2763), .B(n3206), .Z(n5982) );
  HS65_LLS_XOR2X6 U11807 ( .A(n3002), .B(n2754), .Z(n7578) );
  HS65_LLS_XOR2X6 U11808 ( .A(n2645), .B(n187), .Z(n2697) );
  HS65_LLS_XOR2X6 U11809 ( .A(n2673), .B(n140), .Z(n2712) );
  HS65_LL_NAND4ABX3 U11810 ( .A(n5118), .B(n5119), .C(n5120), .D(n5121), .Z(
        n3212) );
  HS65_LL_MX41X7 U11811 ( .D0(n679), .S0(n697), .D1(n685), .S1(n680), .D2(n684), .S2(n677), .D3(n678), .S3(n4638), .Z(n5119) );
  HS65_LL_AOI212X4 U11812 ( .A(n695), .B(n5122), .C(n673), .D(n4854), .E(n5123), .Z(n5121) );
  HS65_LL_MX41X7 U11813 ( .D0(n669), .S0(n701), .D1(n699), .S1(n676), .D2(n702), .S2(n674), .D3(n675), .S3(n688), .Z(n5118) );
  HS65_LLS_XOR2X6 U11814 ( .A(n2803), .B(n572), .Z(n7540) );
  HS65_LLS_XOR2X6 U11815 ( .A(n2819), .B(n230), .Z(n4355) );
  HS65_LLS_XOR2X6 U11816 ( .A(n2811), .B(n2787), .Z(n5948) );
  HS65_LL_NAND4ABX3 U11817 ( .A(n4074), .B(n4075), .C(n4076), .D(n4077), .Z(
        n2674) );
  HS65_LL_MX41X7 U11818 ( .D0(n146), .S0(n169), .D1(n142), .S1(n165), .D2(n147), .S2(n179), .D3(n156), .S3(n166), .Z(n4074) );
  HS65_LL_MX41X7 U11819 ( .D0(n170), .S0(n150), .D1(n180), .S1(n151), .D2(n152), .S2(n168), .D3(n149), .S3(n3040), .Z(n4075) );
  HS65_LL_NOR4ABX2 U11820 ( .A(n3618), .B(n4078), .C(n3030), .D(n3632), .Z(
        n4077) );
  HS65_LL_AOI222X2 U11821 ( .A(n268), .B(n241), .C(n237), .D(n256), .E(n244), 
        .F(n265), .Z(n5313) );
  HS65_LL_AOI222X2 U11822 ( .A(n485), .B(n458), .C(n454), .D(n473), .E(n461), 
        .F(n482), .Z(n5428) );
  HS65_LL_AOI222X2 U11823 ( .A(n82), .B(n57), .C(n58), .D(n74), .E(n55), .F(
        n79), .Z(n6905) );
  HS65_LL_AOI222X2 U11824 ( .A(n694), .B(n669), .C(n673), .D(n686), .E(n670), 
        .F(n695), .Z(n5197) );
  HS65_LL_AOI222X2 U11825 ( .A(n310), .B(n283), .C(n279), .D(n298), .E(n286), 
        .F(n307), .Z(n7020) );
  HS65_LL_AOI222X2 U11826 ( .A(n518), .B(n493), .C(n497), .D(n510), .E(n494), 
        .F(n519), .Z(n6789) );
  HS65_LL_AOI222X2 U11827 ( .A(n283), .B(n304), .C(n286), .D(n310), .E(n297), 
        .F(n284), .Z(n6535) );
  HS65_LL_AOI222X2 U11828 ( .A(n57), .B(n84), .C(n55), .D(n82), .E(n90), .F(
        n54), .Z(n6482) );
  HS65_LL_AOI222X2 U11829 ( .A(n241), .B(n262), .C(n244), .D(n268), .E(n255), 
        .F(n242), .Z(n4889) );
  HS65_LL_AOI222X2 U11830 ( .A(n458), .B(n479), .C(n461), .D(n485), .E(n472), 
        .F(n459), .Z(n4942) );
  HS65_LL_AOI222X2 U11831 ( .A(n493), .B(n515), .C(n494), .D(n518), .E(n523), 
        .F(n495), .Z(n6407) );
  HS65_LL_AOI222X2 U11832 ( .A(n669), .B(n691), .C(n670), .D(n694), .E(n699), 
        .F(n671), .Z(n4814) );
  HS65_LL_NAND3X5 U11833 ( .A(n7816), .B(n7817), .C(n7818), .Z(n7628) );
  HS65_LL_NOR3AX2 U11834 ( .A(n7824), .B(n7825), .C(n7826), .Z(n7817) );
  HS65_LL_NOR3AX2 U11835 ( .A(n7827), .B(n7828), .C(n7829), .Z(n7816) );
  HS65_LL_AOI212X4 U11836 ( .A(n614), .B(n580), .C(n600), .D(n578), .E(n7819), 
        .Z(n7818) );
  HS65_LL_AOI222X2 U11837 ( .A(n218), .B(n188), .C(n215), .D(n197), .E(n219), 
        .F(n202), .Z(n4061) );
  HS65_LL_AOI212X4 U11838 ( .A(n104), .B(n124), .C(n136), .D(n99), .E(n8160), 
        .Z(n8159) );
  HS65_LL_AO12X9 U11839 ( .A(n112), .B(n135), .C(n8161), .Z(n8160) );
  HS65_LL_AOI212X4 U11840 ( .A(n195), .B(n217), .C(n199), .D(n212), .E(n4185), 
        .Z(n4184) );
  HS65_LL_CB4I6X9 U11841 ( .A(n200), .B(n197), .C(n223), .D(n3443), .Z(n4185)
         );
  HS65_LL_AOI222X2 U11842 ( .A(n660), .B(n639), .C(n631), .D(n646), .E(n658), 
        .F(n625), .Z(n4259) );
  HS65_LL_AOI222X2 U11843 ( .A(n102), .B(n131), .C(n120), .D(n105), .E(n129), 
        .F(n113), .Z(n9093) );
  HS65_LL_AOI222X2 U11844 ( .A(n582), .B(n611), .C(n600), .D(n585), .E(n609), 
        .F(n593), .Z(n9035) );
  HS65_LL_AOI222X2 U11845 ( .A(n390), .B(n366), .C(n393), .D(n7963), .E(n363), 
        .F(n396), .Z(n8293) );
  HS65_LL_AOI222X2 U11846 ( .A(n415), .B(n427), .C(n407), .D(n440), .E(n418), 
        .F(n429), .Z(n3810) );
  HS65_LL_AOI222X2 U11847 ( .A(n192), .B(n209), .C(n200), .D(n220), .E(n193), 
        .F(n210), .Z(n3453) );
  HS65_LL_AOI222X2 U11848 ( .A(n147), .B(n172), .C(n165), .D(n155), .E(n148), 
        .F(n173), .Z(n3577) );
  HS65_LL_AOI212X4 U11849 ( .A(n584), .B(n604), .C(n616), .D(n579), .E(n8137), 
        .Z(n8125) );
  HS65_LL_AO12X9 U11850 ( .A(n592), .B(n615), .C(n8138), .Z(n8137) );
  HS65_LL_NAND4ABX3 U11851 ( .A(n4181), .B(n4182), .C(n4183), .D(n4184), .Z(
        n4051) );
  HS65_LL_NAND3AX6 U11852 ( .A(n3488), .B(n3420), .C(n3529), .Z(n4182) );
  HS65_LL_NAND4ABX3 U11853 ( .A(n2954), .B(n3432), .C(n3092), .D(n3510), .Z(
        n4181) );
  HS65_LL_AOI222X2 U11854 ( .A(n188), .B(n224), .C(n219), .D(n203), .E(n209), 
        .F(n201), .Z(n4183) );
  HS65_LL_NAND4ABX3 U11855 ( .A(n8503), .B(n8504), .C(n8505), .D(n8506), .Z(
        n8042) );
  HS65_LL_AOI222X2 U11856 ( .A(n333), .B(n342), .C(n324), .D(n354), .E(n341), 
        .F(n332), .Z(n8505) );
  HS65_LL_NAND4ABX3 U11857 ( .A(n8511), .B(n8512), .C(n8513), .D(n8514), .Z(
        n8504) );
  HS65_LL_AOI212X4 U11858 ( .A(n345), .B(n8507), .C(n349), .D(n8508), .E(n8509), .Z(n8506) );
  HS65_LL_NAND4ABX3 U11859 ( .A(n8200), .B(n8201), .C(n8202), .D(n8203), .Z(
        n7974) );
  HS65_LL_AOI212X4 U11860 ( .A(n384), .B(n8204), .C(n398), .D(n8205), .E(n8206), .Z(n8203) );
  HS65_LL_AOI222X2 U11861 ( .A(n367), .B(n390), .C(n371), .D(n394), .E(n391), 
        .F(n369), .Z(n8202) );
  HS65_LL_NAND4ABX3 U11862 ( .A(n8208), .B(n8209), .C(n8210), .D(n8211), .Z(
        n8201) );
  HS65_LL_NAND4ABX3 U11863 ( .A(n3562), .B(n3563), .C(n3564), .D(n3565), .Z(
        n3227) );
  HS65_LL_NOR3X4 U11864 ( .A(n3566), .B(n3567), .C(n3568), .Z(n3565) );
  HS65_LL_NAND4ABX3 U11865 ( .A(n3569), .B(n3570), .C(n3571), .D(n3572), .Z(
        n3563) );
  HS65_LL_AOI222X2 U11866 ( .A(n142), .B(n172), .C(n166), .D(n3045), .E(n164), 
        .F(n143), .Z(n3564) );
  HS65_LL_NAND4ABX3 U11867 ( .A(n3438), .B(n3439), .C(n3440), .D(n3441), .Z(
        n3071) );
  HS65_LL_NOR3X4 U11868 ( .A(n3442), .B(n3443), .C(n3444), .Z(n3441) );
  HS65_LL_NAND4ABX3 U11869 ( .A(n3445), .B(n3446), .C(n3447), .D(n3448), .Z(
        n3439) );
  HS65_LL_AOI222X2 U11870 ( .A(n209), .B(n188), .C(n221), .D(n2929), .E(n189), 
        .F(n219), .Z(n3440) );
  HS65_LL_NAND4ABX3 U11871 ( .A(n3796), .B(n3797), .C(n3798), .D(n3799), .Z(
        n3356) );
  HS65_LL_AOI222X2 U11872 ( .A(n427), .B(n420), .C(n441), .D(n3195), .E(n422), 
        .F(n442), .Z(n3798) );
  HS65_LL_NOR3AX2 U11873 ( .A(n3800), .B(n3801), .C(n3802), .Z(n3799) );
  HS65_LL_NAND4ABX3 U11874 ( .A(n3803), .B(n2840), .C(n3804), .D(n3805), .Z(
        n3797) );
  HS65_LL_NAND4ABX3 U11875 ( .A(n4082), .B(n4083), .C(n4084), .D(n4085), .Z(
        n3987) );
  HS65_LL_NAND3X5 U11876 ( .A(n3255), .B(n3625), .C(n4096), .Z(n4083) );
  HS65_LL_MX41X7 U11877 ( .D0(n175), .S0(n155), .D1(n153), .S1(n172), .D2(n148), .S2(n163), .D3(n170), .S3(n146), .Z(n4082) );
  HS65_LL_AOI212X4 U11878 ( .A(n166), .B(n3585), .C(n154), .D(n165), .E(n4086), 
        .Z(n4085) );
  HS65_LL_NAND4ABX3 U11879 ( .A(n5646), .B(n5647), .C(n5648), .D(n5649), .Z(
        n5475) );
  HS65_LL_NAND4ABX3 U11880 ( .A(n5024), .B(n5650), .C(n4720), .D(n5003), .Z(
        n5647) );
  HS65_LL_AOI222X2 U11881 ( .A(n11), .B(n40), .C(n24), .D(n45), .E(n39), .F(
        n20), .Z(n5648) );
  HS65_LL_NOR4ABX2 U11882 ( .A(n5066), .B(n4706), .C(n5043), .D(n5098), .Z(
        n5649) );
  HS65_LL_NAND4ABX3 U11883 ( .A(n7238), .B(n7239), .C(n7240), .D(n7241), .Z(
        n7067) );
  HS65_LL_NAND4ABX3 U11884 ( .A(n6617), .B(n7242), .C(n6313), .D(n6596), .Z(
        n7239) );
  HS65_LL_AOI222X2 U11885 ( .A(n533), .B(n562), .C(n546), .D(n567), .E(n561), 
        .F(n542), .Z(n7240) );
  HS65_LL_NOR4ABX2 U11886 ( .A(n6659), .B(n6299), .C(n6636), .D(n6691), .Z(
        n7241) );
  HS65_LL_NAND4ABX3 U11887 ( .A(n8486), .B(n8487), .C(n8488), .D(n8489), .Z(
        n7756) );
  HS65_LL_AOI222X2 U11888 ( .A(n391), .B(n365), .C(n384), .D(n378), .E(n390), 
        .F(n372), .Z(n8488) );
  HS65_LL_NOR4ABX2 U11889 ( .A(n8281), .B(n8107), .C(n8275), .D(n8217), .Z(
        n8489) );
  HS65_LL_MX41X7 U11890 ( .D0(n363), .S0(n395), .D1(n392), .S1(n376), .D2(n377), .S2(n389), .D3(n375), .S3(n398), .Z(n8486) );
  HS65_LL_NAND4ABX3 U11891 ( .A(n5825), .B(n5826), .C(n5827), .D(n5828), .Z(
        n5523) );
  HS65_LL_AOI222X2 U11892 ( .A(n246), .B(n265), .C(n253), .D(n234), .E(n238), 
        .F(n268), .Z(n5827) );
  HS65_LL_NOR4ABX2 U11893 ( .A(n5304), .B(n4919), .C(n5283), .D(n5349), .Z(
        n5828) );
  HS65_LL_NAND4ABX3 U11894 ( .A(n5263), .B(n4930), .C(n5829), .D(n5242), .Z(
        n5826) );
  HS65_LL_NAND4ABX3 U11895 ( .A(n5884), .B(n5885), .C(n5886), .D(n5887), .Z(
        n5545) );
  HS65_LL_AOI222X2 U11896 ( .A(n463), .B(n482), .C(n470), .D(n451), .E(n455), 
        .F(n485), .Z(n5886) );
  HS65_LL_NOR4ABX2 U11897 ( .A(n5419), .B(n4972), .C(n5398), .D(n5464), .Z(
        n5887) );
  HS65_LL_NAND4ABX3 U11898 ( .A(n5378), .B(n4983), .C(n5888), .D(n5357), .Z(
        n5885) );
  HS65_LL_NAND4ABX3 U11899 ( .A(n5676), .B(n5677), .C(n5678), .D(n5679), .Z(
        n5489) );
  HS65_LL_AOI222X2 U11900 ( .A(n668), .B(n695), .C(n700), .D(n679), .E(n675), 
        .F(n694), .Z(n5678) );
  HS65_LL_NOR4ABX2 U11901 ( .A(n5188), .B(n4844), .C(n5166), .D(n5234), .Z(
        n5679) );
  HS65_LL_NAND4ABX3 U11902 ( .A(n5146), .B(n4857), .C(n5680), .D(n5124), .Z(
        n5677) );
  HS65_LL_NAND4ABX3 U11903 ( .A(n7417), .B(n7418), .C(n7419), .D(n7420), .Z(
        n7115) );
  HS65_LL_AOI222X2 U11904 ( .A(n67), .B(n79), .C(n88), .D(n63), .E(n60), .F(
        n82), .Z(n7419) );
  HS65_LL_NOR4ABX2 U11905 ( .A(n6896), .B(n6512), .C(n6875), .D(n6941), .Z(
        n7420) );
  HS65_LL_NAND4ABX3 U11906 ( .A(n6855), .B(n6523), .C(n7421), .D(n6834), .Z(
        n7418) );
  HS65_LL_NAND4ABX3 U11907 ( .A(n7476), .B(n7477), .C(n7478), .D(n7479), .Z(
        n7137) );
  HS65_LL_AOI222X2 U11908 ( .A(n288), .B(n307), .C(n295), .D(n276), .E(n280), 
        .F(n310), .Z(n7478) );
  HS65_LL_NOR4ABX2 U11909 ( .A(n7011), .B(n6565), .C(n6990), .D(n7056), .Z(
        n7479) );
  HS65_LL_NAND4ABX3 U11910 ( .A(n6970), .B(n6576), .C(n7480), .D(n6949), .Z(
        n7477) );
  HS65_LL_NAND4ABX3 U11911 ( .A(n7268), .B(n7269), .C(n7270), .D(n7271), .Z(
        n7081) );
  HS65_LL_AOI222X2 U11912 ( .A(n492), .B(n519), .C(n524), .D(n503), .E(n499), 
        .F(n518), .Z(n7270) );
  HS65_LL_NOR4ABX2 U11913 ( .A(n6780), .B(n6437), .C(n6758), .D(n6826), .Z(
        n7271) );
  HS65_LL_NAND4ABX3 U11914 ( .A(n6738), .B(n6450), .C(n7272), .D(n6716), .Z(
        n7269) );
  HS65_LL_NAND4ABX3 U11915 ( .A(n8070), .B(n8071), .C(n8072), .D(n8073), .Z(
        n7856) );
  HS65_LL_NOR3AX2 U11916 ( .A(n8074), .B(n8075), .C(n8076), .Z(n8073) );
  HS65_LL_AOI222X2 U11917 ( .A(n367), .B(n397), .C(n390), .D(n369), .E(n368), 
        .F(n386), .Z(n8072) );
  HS65_LL_NAND3AX6 U11918 ( .A(n8077), .B(n8078), .C(n8079), .Z(n8071) );
  HS65_LL_NAND4ABX3 U11919 ( .A(n8515), .B(n8516), .C(n8517), .D(n8518), .Z(
        n8315) );
  HS65_LL_NOR3X4 U11920 ( .A(n8519), .B(n8520), .C(n8521), .Z(n8518) );
  HS65_LL_AOI222X2 U11921 ( .A(n342), .B(n322), .C(n355), .D(n8031), .E(n320), 
        .F(n356), .Z(n8517) );
  HS65_LL_NAND4ABX3 U11922 ( .A(n8522), .B(n8523), .C(n8524), .D(n8525), .Z(
        n8516) );
  HS65_LL_NAND4ABX3 U11923 ( .A(n8864), .B(n8865), .C(n8866), .D(n8867), .Z(
        n7774) );
  HS65_LL_NAND4ABX3 U11924 ( .A(n8868), .B(n8323), .C(n8555), .D(n8502), .Z(
        n8865) );
  HS65_LL_AOI222X2 U11925 ( .A(n341), .B(n319), .C(n345), .D(n330), .E(n342), 
        .F(n326), .Z(n8866) );
  HS65_LL_NOR4ABX2 U11926 ( .A(n8586), .B(n8572), .C(n8344), .D(n8606), .Z(
        n8867) );
  HS65_LL_NAND4ABX3 U11927 ( .A(n4059), .B(n4060), .C(n4061), .D(n4062), .Z(
        n3894) );
  HS65_LL_NAND4ABX3 U11928 ( .A(n3121), .B(n3078), .C(n2953), .D(n3091), .Z(
        n4060) );
  HS65_LL_NOR4ABX2 U11929 ( .A(n3521), .B(n3476), .C(n3492), .D(n3512), .Z(
        n4062) );
  HS65_LL_NAND4ABX3 U11930 ( .A(n3442), .B(n3463), .C(n3431), .D(n4063), .Z(
        n4059) );
  HS65_LL_NOR2X6 U11931 ( .A(n168), .B(n163), .Z(n2919) );
  HS65_LL_NOR2X6 U11932 ( .A(n606), .B(n615), .Z(n7618) );
  HS65_LL_NOR2X6 U11933 ( .A(n126), .B(n135), .Z(n7659) );
  HS65_LL_NOR2X6 U11934 ( .A(n515), .B(n508), .Z(n6128) );
  HS65_LL_NOR2X6 U11935 ( .A(n262), .B(n258), .Z(n4587) );
  HS65_LL_NOR2X6 U11936 ( .A(n304), .B(n300), .Z(n6197) );
  HS65_LL_NOR2X6 U11937 ( .A(n84), .B(n73), .Z(n6180) );
  HS65_LL_NOR2X6 U11938 ( .A(n691), .B(n684), .Z(n4535) );
  HS65_LL_NOR2X6 U11939 ( .A(n479), .B(n475), .Z(n4604) );
  HS65_LL_NOR2X6 U11940 ( .A(n438), .B(n443), .Z(n2998) );
  HS65_LL_NOR2X6 U11941 ( .A(n655), .B(n652), .Z(n2973) );
  HS65_LL_NOR2X6 U11942 ( .A(n214), .B(n218), .Z(n2861) );
  HS65_LL_NOR2X6 U11943 ( .A(n558), .B(n551), .Z(n6072) );
  HS65_LL_NOR2X6 U11944 ( .A(n36), .B(n29), .Z(n4479) );
  HS65_LL_NOR2X6 U11945 ( .A(n397), .B(n395), .Z(n7852) );
  HS65_LL_NOR2X6 U11946 ( .A(n352), .B(n353), .Z(n7953) );
  HS65_LL_NAND4ABX3 U11947 ( .A(n5712), .B(n5713), .C(n5714), .D(n5715), .Z(
        n5645) );
  HS65_LL_NAND3AX6 U11948 ( .A(n5022), .B(n5065), .C(n5004), .Z(n5713) );
  HS65_LL_AOI222X2 U11949 ( .A(n9), .B(n45), .C(n20), .D(n30), .E(n39), .F(n19), .Z(n5714) );
  HS65_LL_NAND4ABX3 U11950 ( .A(n4564), .B(n4707), .C(n5096), .D(n5041), .Z(
        n5712) );
  HS65_LL_NAND4ABX3 U11951 ( .A(n7304), .B(n7305), .C(n7306), .D(n7307), .Z(
        n7237) );
  HS65_LL_NAND3AX6 U11952 ( .A(n6615), .B(n6658), .C(n6597), .Z(n7305) );
  HS65_LL_AOI222X2 U11953 ( .A(n531), .B(n567), .C(n542), .D(n552), .E(n561), 
        .F(n541), .Z(n7306) );
  HS65_LL_NAND4ABX3 U11954 ( .A(n6157), .B(n6300), .C(n6689), .D(n6634), .Z(
        n7304) );
  HS65_LL_NAND4ABX3 U11955 ( .A(n7900), .B(n7901), .C(n7902), .D(n7903), .Z(
        n7718) );
  HS65_LL_AOI222X2 U11956 ( .A(n104), .B(n120), .C(n136), .D(n113), .E(n112), 
        .F(n129), .Z(n7902) );
  HS65_LL_NAND3X5 U11957 ( .A(n7907), .B(n7908), .C(n7909), .Z(n7901) );
  HS65_LL_NAND4ABX3 U11958 ( .A(n7910), .B(n7911), .C(n7912), .D(n7913), .Z(
        n7900) );
  HS65_LL_NAND4ABX3 U11959 ( .A(n7801), .B(n7802), .C(n7803), .D(n7804), .Z(
        n7680) );
  HS65_LL_AOI222X2 U11960 ( .A(n584), .B(n600), .C(n616), .D(n593), .E(n592), 
        .F(n609), .Z(n7803) );
  HS65_LL_NAND3X5 U11961 ( .A(n7809), .B(n7810), .C(n7811), .Z(n7802) );
  HS65_LL_NAND4ABX3 U11962 ( .A(n7812), .B(n7813), .C(n7814), .D(n7815), .Z(
        n7801) );
  HS65_LL_NAND3X5 U11963 ( .A(n5618), .B(n5619), .C(n5620), .Z(n4513) );
  HS65_LL_AND3X9 U11964 ( .A(n4971), .B(n5404), .C(n5418), .Z(n5619) );
  HS65_LL_NOR3X4 U11965 ( .A(n5624), .B(n5384), .C(n5465), .Z(n5618) );
  HS65_LL_AOI212X4 U11966 ( .A(n460), .B(n474), .C(n470), .D(n461), .E(n5621), 
        .Z(n5620) );
  HS65_LL_NAND3X5 U11967 ( .A(n5593), .B(n5594), .C(n5595), .Z(n4452) );
  HS65_LL_AND3X9 U11968 ( .A(n4918), .B(n5289), .C(n5303), .Z(n5594) );
  HS65_LL_NOR3X4 U11969 ( .A(n5599), .B(n5269), .C(n5350), .Z(n5593) );
  HS65_LL_AOI212X4 U11970 ( .A(n243), .B(n257), .C(n253), .D(n244), .E(n5596), 
        .Z(n5595) );
  HS65_LL_NAND3X5 U11971 ( .A(n7210), .B(n7211), .C(n7212), .Z(n6106) );
  HS65_LL_AND3X9 U11972 ( .A(n6564), .B(n6996), .C(n7010), .Z(n7211) );
  HS65_LL_NOR3X4 U11973 ( .A(n7216), .B(n6976), .C(n7057), .Z(n7210) );
  HS65_LL_AOI212X4 U11974 ( .A(n285), .B(n299), .C(n295), .D(n286), .E(n7213), 
        .Z(n7212) );
  HS65_LL_NAND3X5 U11975 ( .A(n5767), .B(n5768), .C(n5769), .Z(n5569) );
  HS65_LL_AND3X9 U11976 ( .A(n4843), .B(n5173), .C(n5187), .Z(n5768) );
  HS65_LL_NOR3X4 U11977 ( .A(n5773), .B(n5152), .C(n5235), .Z(n5767) );
  HS65_LL_AOI212X4 U11978 ( .A(n672), .B(n688), .C(n700), .D(n670), .E(n5770), 
        .Z(n5769) );
  HS65_LL_NAND3X5 U11979 ( .A(n7359), .B(n7360), .C(n7361), .Z(n7161) );
  HS65_LL_AND3X9 U11980 ( .A(n6436), .B(n6765), .C(n6779), .Z(n7360) );
  HS65_LL_NOR3X4 U11981 ( .A(n7365), .B(n6744), .C(n6827), .Z(n7359) );
  HS65_LL_AOI212X4 U11982 ( .A(n496), .B(n512), .C(n524), .D(n494), .E(n7362), 
        .Z(n7361) );
  HS65_LL_NAND3X5 U11983 ( .A(n4112), .B(n4113), .C(n4114), .Z(n3986) );
  HS65_LL_NOR3X4 U11984 ( .A(n3630), .B(n3645), .C(n3616), .Z(n4113) );
  HS65_LL_NOR3X4 U11985 ( .A(n4118), .B(n3245), .C(n3556), .Z(n4112) );
  HS65_LL_AOI212X4 U11986 ( .A(n166), .B(n149), .C(n148), .D(n178), .E(n4115), 
        .Z(n4114) );
  HS65_LL_NAND3X5 U11987 ( .A(n5705), .B(n5706), .C(n5707), .Z(n5505) );
  HS65_LL_NOR3AX2 U11988 ( .A(n4705), .B(n5050), .C(n5068), .Z(n5706) );
  HS65_LL_NOR3AX2 U11989 ( .A(n5031), .B(n5711), .C(n5099), .Z(n5705) );
  HS65_LL_AOI212X4 U11990 ( .A(n17), .B(n33), .C(n15), .D(n45), .E(n5708), .Z(
        n5707) );
  HS65_LL_NAND3X5 U11991 ( .A(n7297), .B(n7298), .C(n7299), .Z(n7097) );
  HS65_LL_NOR3AX2 U11992 ( .A(n6298), .B(n6643), .C(n6661), .Z(n7298) );
  HS65_LL_NOR3AX2 U11993 ( .A(n6624), .B(n7303), .C(n6692), .Z(n7297) );
  HS65_LL_AOI212X4 U11994 ( .A(n539), .B(n555), .C(n537), .D(n567), .E(n7300), 
        .Z(n7299) );
  HS65_LL_NAND4ABX3 U11995 ( .A(n6747), .B(n6748), .C(n6749), .D(n6750), .Z(
        n6427) );
  HS65_LL_NAND3X5 U11996 ( .A(n6759), .B(n6760), .C(n6761), .Z(n6748) );
  HS65_LL_NOR4ABX2 U11997 ( .A(n6751), .B(n6752), .C(n6753), .D(n6754), .Z(
        n6750) );
  HS65_LL_NAND4ABX3 U11998 ( .A(n6763), .B(n6764), .C(n6765), .D(n6766), .Z(
        n6747) );
  HS65_LL_NAND4ABX3 U11999 ( .A(n5155), .B(n5156), .C(n5157), .D(n5158), .Z(
        n4834) );
  HS65_LL_NAND3X5 U12000 ( .A(n5167), .B(n5168), .C(n5169), .Z(n5156) );
  HS65_LL_NOR4ABX2 U12001 ( .A(n5159), .B(n5160), .C(n5161), .D(n5162), .Z(
        n5158) );
  HS65_LL_NAND4ABX3 U12002 ( .A(n5171), .B(n5172), .C(n5173), .D(n5174), .Z(
        n5155) );
  HS65_LL_NAND4ABX3 U12003 ( .A(n5387), .B(n5388), .C(n5389), .D(n5390), .Z(
        n4962) );
  HS65_LL_NAND3X5 U12004 ( .A(n5399), .B(n5400), .C(n5401), .Z(n5388) );
  HS65_LL_NOR4ABX2 U12005 ( .A(n5391), .B(n5392), .C(n5393), .D(n5394), .Z(
        n5390) );
  HS65_LL_NAND4ABX3 U12006 ( .A(n5402), .B(n5403), .C(n5404), .D(n5405), .Z(
        n5387) );
  HS65_LL_NAND4ABX3 U12007 ( .A(n8560), .B(n8561), .C(n8562), .D(n8563), .Z(
        n8326) );
  HS65_LL_NAND3AX6 U12008 ( .A(n7764), .B(n8572), .C(n8573), .Z(n8561) );
  HS65_LL_NOR4ABX2 U12009 ( .A(n8564), .B(n8565), .C(n8566), .D(n8567), .Z(
        n8563) );
  HS65_LL_NOR4ABX2 U12010 ( .A(n8568), .B(n8569), .C(n8570), .D(n8571), .Z(
        n8562) );
  HS65_LL_NAND4ABX3 U12011 ( .A(n6626), .B(n6627), .C(n6628), .D(n6629), .Z(
        n6289) );
  HS65_LL_NOR4ABX2 U12012 ( .A(n6634), .B(n6635), .C(n6636), .D(n6637), .Z(
        n6628) );
  HS65_LL_NAND3X5 U12013 ( .A(n6638), .B(n6639), .C(n6640), .Z(n6627) );
  HS65_LL_NOR4ABX2 U12014 ( .A(n6630), .B(n6631), .C(n6632), .D(n6633), .Z(
        n6629) );
  HS65_LL_NAND4ABX3 U12015 ( .A(n5033), .B(n5034), .C(n5035), .D(n5036), .Z(
        n4696) );
  HS65_LL_NOR4ABX2 U12016 ( .A(n5041), .B(n5042), .C(n5043), .D(n5044), .Z(
        n5035) );
  HS65_LL_NAND3X5 U12017 ( .A(n5045), .B(n5046), .C(n5047), .Z(n5034) );
  HS65_LL_NOR4ABX2 U12018 ( .A(n5037), .B(n5038), .C(n5039), .D(n5040), .Z(
        n5036) );
  HS65_LL_NAND4ABX3 U12019 ( .A(n3228), .B(n3229), .C(n3230), .D(n3231), .Z(
        n3020) );
  HS65_LL_NAND4ABX3 U12020 ( .A(n3259), .B(n3260), .C(n3261), .D(n3262), .Z(
        n3229) );
  HS65_LL_NOR4ABX2 U12021 ( .A(n3232), .B(n3233), .C(n3234), .D(n3235), .Z(
        n3231) );
  HS65_LL_MX41X7 U12022 ( .D0(n168), .S0(n146), .D1(n175), .S1(n143), .D2(n156), .S2(n177), .D3(n152), .S3(n172), .Z(n3228) );
  HS65_LL_OAI31X5 U12023 ( .A(n606), .B(n612), .C(n614), .D(n582), .Z(n8381)
         );
  HS65_LL_OAI31X5 U12024 ( .A(n126), .B(n132), .C(n134), .D(n102), .Z(n8433)
         );
  HS65_LL_NAND4ABX3 U12025 ( .A(n8316), .B(n8317), .C(n8318), .D(n8319), .Z(
        n8043) );
  HS65_LL_NAND4ABX3 U12026 ( .A(n8345), .B(n8346), .C(n8347), .D(n8348), .Z(
        n8317) );
  HS65_LL_MX41X7 U12027 ( .D0(n317), .S0(n352), .D1(n343), .S1(n320), .D2(n323), .S2(n347), .D3(n342), .S3(n327), .Z(n8316) );
  HS65_LL_NOR4ABX2 U12028 ( .A(n8320), .B(n8321), .C(n8322), .D(n8323), .Z(
        n8319) );
  HS65_LL_NAND4ABX3 U12029 ( .A(n3072), .B(n3073), .C(n3074), .D(n3075), .Z(
        n2944) );
  HS65_LL_NAND4ABX3 U12030 ( .A(n3103), .B(n3104), .C(n3105), .D(n3106), .Z(
        n3073) );
  HS65_LL_NOR4ABX2 U12031 ( .A(n3076), .B(n3077), .C(n3078), .D(n3079), .Z(
        n3075) );
  HS65_LL_MX41X7 U12032 ( .D0(n191), .S0(n214), .D1(n189), .S1(n211), .D2(n201), .S2(n223), .D3(n197), .S3(n209), .Z(n3072) );
  HS65_LL_NAND4ABX3 U12033 ( .A(n8084), .B(n8085), .C(n8086), .D(n8087), .Z(
        n7975) );
  HS65_LL_NAND4ABX3 U12034 ( .A(n8112), .B(n8113), .C(n8114), .D(n8115), .Z(
        n8085) );
  HS65_LL_MX41X7 U12035 ( .D0(n362), .S0(n397), .D1(n392), .S1(n363), .D2(n373), .S2(n386), .D3(n390), .S3(n375), .Z(n8084) );
  HS65_LL_NOR4ABX2 U12036 ( .A(n8088), .B(n8089), .C(n8090), .D(n8091), .Z(
        n8087) );
  HS65_LL_OAI31X5 U12037 ( .A(n343), .B(n352), .C(n355), .D(n319), .Z(n8320)
         );
  HS65_LL_NAND4ABX3 U12038 ( .A(n8833), .B(n8834), .C(n8835), .D(n8836), .Z(
        n8162) );
  HS65_LL_AOI222X2 U12039 ( .A(n129), .B(n99), .C(n111), .D(n137), .E(n98), 
        .F(n131), .Z(n8835) );
  HS65_LL_AOI212X4 U12040 ( .A(n120), .B(n7722), .C(n124), .D(n8837), .E(n8838), .Z(n8836) );
  HS65_LL_NAND4ABX3 U12041 ( .A(n8839), .B(n8840), .C(n7890), .D(n8841), .Z(
        n8834) );
  HS65_LL_OAI31X5 U12042 ( .A(n211), .B(n214), .C(n221), .D(n190), .Z(n3076)
         );
  HS65_LL_OAI31X5 U12043 ( .A(n392), .B(n397), .C(n393), .D(n365), .Z(n8088)
         );
  HS65_LL_OAI31X5 U12044 ( .A(n264), .B(n257), .C(n262), .D(n246), .Z(n4904)
         );
  HS65_LL_OAI31X5 U12045 ( .A(n481), .B(n474), .C(n479), .D(n463), .Z(n4957)
         );
  HS65_LL_OAI31X5 U12046 ( .A(n306), .B(n299), .C(n304), .D(n288), .Z(n6550)
         );
  HS65_LL_OAI31X5 U12047 ( .A(n78), .B(n76), .C(n84), .D(n67), .Z(n6497) );
  HS65_LL_OAI31X5 U12048 ( .A(n521), .B(n512), .C(n515), .D(n492), .Z(n6422)
         );
  HS65_LL_OAI31X5 U12049 ( .A(n697), .B(n688), .C(n691), .D(n668), .Z(n4829)
         );
  HS65_LL_OAI31X5 U12050 ( .A(n661), .B(n655), .C(n650), .D(n639), .Z(n3307)
         );
  HS65_LL_OAI31X5 U12051 ( .A(n430), .B(n438), .C(n441), .D(n421), .Z(n3361)
         );
  HS65_LL_NAND4ABX3 U12052 ( .A(n3021), .B(n3022), .C(n3023), .D(n3024), .Z(
        n2909) );
  HS65_LL_NOR3AX2 U12053 ( .A(n3029), .B(n3030), .C(n3031), .Z(n3023) );
  HS65_LL_NOR4ABX2 U12054 ( .A(n3025), .B(n3026), .C(n3027), .D(n3028), .Z(
        n3024) );
  HS65_LL_NAND3AX6 U12055 ( .A(n3037), .B(n3038), .C(n3039), .Z(n3021) );
  HS65_LL_OAI31X5 U12056 ( .A(n175), .B(n166), .C(n168), .D(n145), .Z(n3232)
         );
  HS65_LL_OAI31X5 U12057 ( .A(n42), .B(n33), .C(n36), .D(n11), .Z(n4691) );
  HS65_LL_OAI31X5 U12058 ( .A(n564), .B(n555), .C(n558), .D(n533), .Z(n6284)
         );
  HS65_LL_NOR2X6 U12059 ( .A(n780), .B(n785), .Z(n1950) );
  HS65_LL_NOR2X6 U12060 ( .A(n862), .B(n867), .Z(n1198) );
  HS65_LL_NOR3X4 U12061 ( .A(n3609), .B(n3027), .C(n3644), .Z(n4096) );
  HS65_LL_NOR3X4 U12062 ( .A(n7857), .B(n8092), .C(n8093), .Z(n8086) );
  HS65_LL_NOR2X6 U12063 ( .A(n903), .B(n908), .Z(n2326) );
  HS65_LL_NOR2X6 U12064 ( .A(n821), .B(n826), .Z(n1574) );
  HS65_LL_NOR3X4 U12065 ( .A(n7998), .B(n8386), .C(n8387), .Z(n8379) );
  HS65_LL_NOR3X4 U12066 ( .A(n8011), .B(n8438), .C(n8439), .Z(n8431) );
  HS65_LL_NOR2X6 U12067 ( .A(n177), .B(n170), .Z(n3041) );
  HS65_LL_NOR2X6 U12068 ( .A(n44), .B(n37), .Z(n4565) );
  HS65_LL_NOR2X6 U12069 ( .A(n566), .B(n559), .Z(n6158) );
  HS65_LL_NAND4ABX3 U12070 ( .A(n4297), .B(n4298), .C(n4299), .D(n4300), .Z(
        n3960) );
  HS65_LL_NAND4ABX3 U12071 ( .A(n3402), .B(n3363), .C(n3180), .D(n3376), .Z(
        n4298) );
  HS65_LL_AOI222X2 U12072 ( .A(n443), .B(n420), .C(n437), .D(n411), .E(n442), 
        .F(n408), .Z(n4299) );
  HS65_LL_NAND4ABX3 U12073 ( .A(n3801), .B(n3820), .C(n3789), .D(n4301), .Z(
        n4297) );
  HS65_LL_NOR3X4 U12074 ( .A(n3237), .B(n3238), .C(n2910), .Z(n3230) );
  HS65_LL_NOR3X4 U12075 ( .A(n3081), .B(n3082), .C(n2867), .Z(n3074) );
  HS65_LL_NOR2X6 U12076 ( .A(n599), .B(n615), .Z(n8719) );
  HS65_LL_NOR2X6 U12077 ( .A(n119), .B(n135), .Z(n8809) );
  HS65_LL_NOR2X6 U12078 ( .A(n472), .B(n475), .Z(n5559) );
  HS65_LL_NOR2X6 U12079 ( .A(n255), .B(n258), .Z(n5537) );
  HS65_LL_NOR2X6 U12080 ( .A(n699), .B(n684), .Z(n5494) );
  HS65_LL_NOR2X6 U12081 ( .A(n297), .B(n300), .Z(n7151) );
  HS65_LL_NOR2X6 U12082 ( .A(n523), .B(n508), .Z(n7086) );
  HS65_LL_NOR2X6 U12083 ( .A(n90), .B(n73), .Z(n7129) );
  HS65_LL_NOR2X6 U12084 ( .A(n342), .B(n340), .Z(n8542) );
  HS65_LL_NOR2X6 U12085 ( .A(n209), .B(n212), .Z(n3477) );
  HS65_LL_NOR2X6 U12086 ( .A(n223), .B(n218), .Z(n3890) );
  HS65_LL_NOR2X6 U12087 ( .A(n44), .B(n29), .Z(n5470) );
  HS65_LL_NOR2X6 U12088 ( .A(n566), .B(n551), .Z(n7062) );
  HS65_LL_NAND4ABX3 U12089 ( .A(n5689), .B(n5690), .C(n5691), .D(n5692), .Z(
        n5491) );
  HS65_LL_AOI222X2 U12090 ( .A(n665), .B(n684), .C(n678), .D(n692), .E(n676), 
        .F(n685), .Z(n5691) );
  HS65_LL_NAND4ABX3 U12091 ( .A(n4632), .B(n5143), .C(n5229), .D(n4839), .Z(
        n5690) );
  HS65_LL_NOR4ABX2 U12092 ( .A(n5194), .B(n5183), .C(n5203), .D(n5162), .Z(
        n5692) );
  HS65_LL_NAND4ABX3 U12093 ( .A(n7281), .B(n7282), .C(n7283), .D(n7284), .Z(
        n7083) );
  HS65_LL_AOI222X2 U12094 ( .A(n489), .B(n508), .C(n502), .D(n516), .E(n500), 
        .F(n509), .Z(n7283) );
  HS65_LL_NAND4ABX3 U12095 ( .A(n6225), .B(n6735), .C(n6821), .D(n6432), .Z(
        n7282) );
  HS65_LL_NOR4ABX2 U12096 ( .A(n6786), .B(n6775), .C(n6795), .D(n6754), .Z(
        n7284) );
  HS65_LL_NOR2X6 U12097 ( .A(n694), .B(n696), .Z(n5134) );
  HS65_LL_NOR2X6 U12098 ( .A(n518), .B(n520), .Z(n6726) );
  HS65_LL_NOR2X6 U12099 ( .A(n310), .B(n309), .Z(n6959) );
  HS65_LL_NOR2X6 U12100 ( .A(n82), .B(n81), .Z(n6844) );
  HS65_LL_NOR2X6 U12101 ( .A(n268), .B(n267), .Z(n5252) );
  HS65_LL_NOR2X6 U12102 ( .A(n485), .B(n484), .Z(n5367) );
  HS65_LL_NOR2X6 U12103 ( .A(n39), .B(n41), .Z(n5012) );
  HS65_LL_NOR2X6 U12104 ( .A(n561), .B(n563), .Z(n6605) );
  HS65_LL_NOR2X6 U12105 ( .A(n427), .B(n428), .Z(n3832) );
  HS65_LL_NOR2X6 U12106 ( .A(n609), .B(n610), .Z(n8677) );
  HS65_LL_NOR2X6 U12107 ( .A(n129), .B(n130), .Z(n8767) );
  HS65_LL_NOR2X6 U12108 ( .A(n386), .B(n395), .Z(n8481) );
  HS65_LL_NOR2X6 U12109 ( .A(n172), .B(n174), .Z(n3601) );
  HS65_LL_NOR4ABX2 U12110 ( .A(n4066), .B(n4067), .C(n4068), .D(n4069), .Z(
        n3892) );
  HS65_LL_NAND4ABX3 U12111 ( .A(n3079), .B(n3434), .C(n4070), .D(n3421), .Z(
        n4069) );
  HS65_LL_MX41X7 U12112 ( .D0(n189), .S0(n218), .D1(n211), .S1(n199), .D2(n212), .S2(n196), .D3(n197), .S3(n213), .Z(n4068) );
  HS65_LL_AOI222X2 U12113 ( .A(n210), .B(n190), .C(n198), .D(n224), .E(n209), 
        .F(n203), .Z(n4066) );
  HS65_LL_NOR4ABX2 U12114 ( .A(n9093), .B(n9094), .C(n9095), .D(n9096), .Z(
        n7716) );
  HS65_LL_NAND4ABX3 U12115 ( .A(n8779), .B(n8435), .C(n9097), .D(n8758), .Z(
        n9096) );
  HS65_LL_MX41X7 U12116 ( .D0(n135), .S0(n103), .D1(n107), .S1(n132), .D2(n108), .S2(n130), .D3(n124), .S3(n106), .Z(n9095) );
  HS65_LL_NOR4ABX2 U12117 ( .A(n8803), .B(n8446), .C(n8793), .D(n8821), .Z(
        n9094) );
  HS65_LL_NOR4ABX2 U12118 ( .A(n9035), .B(n9036), .C(n9037), .D(n9038), .Z(
        n7678) );
  HS65_LL_NAND4ABX3 U12119 ( .A(n8689), .B(n8383), .C(n9039), .D(n8668), .Z(
        n9038) );
  HS65_LL_MX41X7 U12120 ( .D0(n615), .S0(n583), .D1(n587), .S1(n612), .D2(n588), .S2(n610), .D3(n604), .S3(n586), .Z(n9037) );
  HS65_LL_NOR4ABX2 U12121 ( .A(n8713), .B(n8394), .C(n8703), .D(n8731), .Z(
        n9036) );
  HS65_LL_NAND4ABX3 U12122 ( .A(n8212), .B(n8213), .C(n8214), .D(n8215), .Z(
        n8093) );
  HS65_LL_NOR3AX2 U12123 ( .A(n8216), .B(n8217), .C(n8218), .Z(n8215) );
  HS65_LL_NAND4ABX3 U12124 ( .A(n8224), .B(n8225), .C(n8226), .D(n8227), .Z(
        n8212) );
  HS65_LL_MX41X7 U12125 ( .D0(n369), .S0(n389), .D1(n373), .S1(n384), .D2(n395), .S2(n370), .D3(n371), .S3(n398), .Z(n8213) );
  HS65_LL_NOR3X4 U12126 ( .A(n8256), .B(n7983), .C(n8276), .Z(n8943) );
  HS65_LL_NOR3X4 U12127 ( .A(n8558), .B(n8051), .C(n8576), .Z(n8883) );
  HS65_LL_NAND2X7 U12128 ( .A(n23), .B(n45), .Z(n5004) );
  HS65_LL_NAND2X7 U12129 ( .A(n545), .B(n567), .Z(n6597) );
  HS65_LL_NAND4ABX3 U12130 ( .A(n3620), .B(n3621), .C(n3622), .D(n3623), .Z(
        n3238) );
  HS65_LL_NOR4ABX2 U12131 ( .A(n3628), .B(n3629), .C(n3630), .D(n3631), .Z(
        n3622) );
  HS65_LL_NOR4ABX2 U12132 ( .A(n3624), .B(n3625), .C(n3626), .D(n3627), .Z(
        n3623) );
  HS65_LL_NAND3AX6 U12133 ( .A(n3632), .B(n3633), .C(n3634), .Z(n3621) );
  HS65_LL_NOR4ABX2 U12134 ( .A(n4259), .B(n4260), .C(n4261), .D(n4262), .Z(
        n3938) );
  HS65_LL_NAND4ABX3 U12135 ( .A(n3310), .B(n3677), .C(n4263), .D(n3664), .Z(
        n4262) );
  HS65_LL_MX41X7 U12136 ( .D0(n640), .S0(n652), .D1(n661), .S1(n630), .D2(n659), .S2(n628), .D3(n629), .S3(n656), .Z(n4261) );
  HS65_LL_NOR4ABX2 U12137 ( .A(n3328), .B(n3759), .C(n3733), .D(n3752), .Z(
        n4260) );
  HS65_LL_NOR4ABX2 U12138 ( .A(n4318), .B(n4319), .C(n4320), .D(n4321), .Z(
        n3958) );
  HS65_LL_NAND4ABX3 U12139 ( .A(n3364), .B(n3792), .C(n4322), .D(n3777), .Z(
        n4321) );
  HS65_LL_MX41X7 U12140 ( .D0(n422), .S0(n443), .D1(n430), .S1(n412), .D2(n428), .S2(n409), .D3(n411), .S3(n439), .Z(n4320) );
  HS65_LL_AOI222X2 U12141 ( .A(n429), .B(n421), .C(n413), .D(n433), .E(n427), 
        .F(n406), .Z(n4318) );
  HS65_LL_NAND3X5 U12142 ( .A(n8720), .B(n8721), .C(n8722), .Z(n8387) );
  HS65_LL_NOR4ABX2 U12143 ( .A(n8727), .B(n7688), .C(n8728), .D(n7793), .Z(
        n8721) );
  HS65_LL_NOR4ABX2 U12144 ( .A(n8729), .B(n7827), .C(n8730), .D(n8731), .Z(
        n8720) );
  HS65_LL_NOR4ABX2 U12145 ( .A(n7814), .B(n8723), .C(n8724), .D(n8725), .Z(
        n8722) );
  HS65_LL_NAND2X7 U12146 ( .A(n175), .B(n147), .Z(n3584) );
  HS65_LL_NAND2X7 U12147 ( .A(n152), .B(n166), .Z(n3558) );
  HS65_LL_NAND2X7 U12148 ( .A(n148), .B(n169), .Z(n3639) );
  HS65_LL_NAND2X7 U12149 ( .A(n580), .B(n616), .Z(n8398) );
  HS65_LL_NAND2X7 U12150 ( .A(n179), .B(n157), .Z(n3596) );
  HS65_LL_NOR2X6 U12151 ( .A(n768), .B(n770), .Z(n1907) );
  HS65_LL_NOR2X6 U12152 ( .A(n891), .B(n893), .Z(n2283) );
  HS65_LL_NOR2X6 U12153 ( .A(n386), .B(n399), .Z(n7959) );
  HS65_LL_NOR2X6 U12154 ( .A(n347), .B(n350), .Z(n8027) );
  HS65_LL_NOR2X6 U12155 ( .A(n255), .B(n261), .Z(n4726) );
  HS65_LL_NOR2X6 U12156 ( .A(n472), .B(n478), .Z(n4788) );
  HS65_LL_NOR2X6 U12157 ( .A(n297), .B(n303), .Z(n6381) );
  HS65_LL_NOR2X6 U12158 ( .A(n90), .B(n85), .Z(n6342) );
  HS65_LL_NOR2X6 U12159 ( .A(n523), .B(n516), .Z(n6235) );
  HS65_LL_NOR2X6 U12160 ( .A(n699), .B(n692), .Z(n4642) );
  HS65_LL_NAND2X7 U12161 ( .A(n332), .B(n351), .Z(n8568) );
  HS65_LL_NOR2X6 U12162 ( .A(n809), .B(n811), .Z(n1531) );
  HS65_LL_NOR2X6 U12163 ( .A(n599), .B(n605), .Z(n7637) );
  HS65_LL_NOR2X6 U12164 ( .A(n119), .B(n125), .Z(n7658) );
  HS65_LL_NOR2X6 U12165 ( .A(n435), .B(n437), .Z(n3191) );
  HS65_LL_NOR2X6 U12166 ( .A(n223), .B(n215), .Z(n2925) );
  HS65_LL_NAND2X7 U12167 ( .A(n499), .B(n524), .Z(n6452) );
  HS65_LL_NAND2X7 U12168 ( .A(n675), .B(n700), .Z(n4859) );
  HS65_LL_NAND2X7 U12169 ( .A(n629), .B(n646), .Z(n3663) );
  HS65_LL_NAND4ABX3 U12170 ( .A(n3422), .B(n3423), .C(n3424), .D(n3425), .Z(
        n3081) );
  HS65_LL_NOR4ABX2 U12171 ( .A(n3426), .B(n3427), .C(n3428), .D(n3429), .Z(
        n3425) );
  HS65_LL_NAND3AX6 U12172 ( .A(n3434), .B(n3435), .C(n3436), .Z(n3422) );
  HS65_LL_NOR4ABX2 U12173 ( .A(n3430), .B(n3431), .C(n3432), .D(n3433), .Z(
        n3424) );
  HS65_LL_NOR2X6 U12174 ( .A(n648), .B(n654), .Z(n3127) );
  HS65_LL_CBI4I6X5 U12175 ( .A(n163), .B(n169), .C(n158), .D(n3566), .Z(n3993)
         );
  HS65_LL_NOR2X6 U12176 ( .A(n804), .B(n799), .Z(n1525) );
  HS65_LL_NAND4ABX3 U12177 ( .A(n4097), .B(n4098), .C(n4099), .D(n4100), .Z(
        n3907) );
  HS65_LL_AOI222X2 U12178 ( .A(n145), .B(n173), .C(n153), .D(n178), .E(n158), 
        .F(n172), .Z(n4099) );
  HS65_LL_NOR4ABX2 U12179 ( .A(n3248), .B(n3646), .C(n3617), .D(n3626), .Z(
        n4100) );
  HS65_LL_NAND4ABX3 U12180 ( .A(n3235), .B(n3555), .C(n4101), .D(n3545), .Z(
        n4098) );
  HS65_LL_NAND4ABX3 U12181 ( .A(n3546), .B(n3547), .C(n3548), .D(n3549), .Z(
        n3237) );
  HS65_LL_NOR4X4 U12182 ( .A(n3554), .B(n3555), .C(n3556), .D(n3557), .Z(n3548) );
  HS65_LL_NOR4ABX2 U12183 ( .A(n3550), .B(n3551), .C(n3552), .D(n3553), .Z(
        n3549) );
  HS65_LL_NAND3X5 U12184 ( .A(n3558), .B(n3559), .C(n3560), .Z(n3546) );
  HS65_LL_NAND2X7 U12185 ( .A(n673), .B(n694), .Z(n5180) );
  HS65_LL_NAND2X7 U12186 ( .A(n497), .B(n518), .Z(n6772) );
  HS65_LL_NAND2X7 U12187 ( .A(n677), .B(n691), .Z(n5216) );
  HS65_LL_NAND2X7 U12188 ( .A(n146), .B(n175), .Z(n3583) );
  HS65_LL_NAND2X7 U12189 ( .A(n106), .B(n127), .Z(n7906) );
  HS65_LL_NAND2X7 U12190 ( .A(n586), .B(n607), .Z(n7808) );
  HS65_LL_NAND2X7 U12191 ( .A(n170), .B(n147), .Z(n3261) );
  HS65_LL_NAND2X7 U12192 ( .A(n154), .B(n170), .Z(n3559) );
  HS65_LL_NAND2X7 U12193 ( .A(n157), .B(n169), .Z(n3051) );
  HS65_LL_NAND4ABX3 U12194 ( .A(n4119), .B(n4120), .C(n4121), .D(n4122), .Z(
        n4088) );
  HS65_LL_AOI222X2 U12195 ( .A(n145), .B(n178), .C(n175), .D(n153), .E(n180), 
        .F(n143), .Z(n4121) );
  HS65_LL_NAND4ABX3 U12196 ( .A(n3568), .B(n3561), .C(n4123), .D(n3583), .Z(
        n4119) );
  HS65_LL_NAND4ABX3 U12197 ( .A(n3249), .B(n3273), .C(n3261), .D(n3025), .Z(
        n4120) );
  HS65_LL_NAND2X7 U12198 ( .A(n56), .B(n74), .Z(n6919) );
  HS65_LL_NAND2X7 U12199 ( .A(n243), .B(n256), .Z(n5327) );
  HS65_LL_NAND2X7 U12200 ( .A(n672), .B(n686), .Z(n5211) );
  HS65_LL_NAND2X7 U12201 ( .A(n496), .B(n510), .Z(n6803) );
  HS65_LL_NOR4ABX2 U12202 ( .A(n5487), .B(n5488), .C(n5489), .D(n5490), .Z(
        n5486) );
  HS65_LL_AOI212X4 U12203 ( .A(n700), .B(n669), .C(n666), .D(n701), .E(n5491), 
        .Z(n5488) );
  HS65_LL_NOR4ABX2 U12204 ( .A(n7079), .B(n7080), .C(n7081), .D(n7082), .Z(
        n7078) );
  HS65_LL_AOI212X4 U12205 ( .A(n524), .B(n493), .C(n490), .D(n525), .E(n7083), 
        .Z(n7080) );
  HS65_LL_NOR2X6 U12206 ( .A(n11), .B(n21), .Z(n4660) );
  HS65_LL_NOR2X6 U12207 ( .A(n533), .B(n543), .Z(n6253) );
  HS65_LL_NAND2X7 U12208 ( .A(n192), .B(n216), .Z(n3435) );
  HS65_LL_NOR2X6 U12209 ( .A(n190), .B(n202), .Z(n3060) );
  HS65_LL_NOR2X6 U12210 ( .A(n639), .B(n627), .Z(n3292) );
  HS65_LL_NOR2X6 U12211 ( .A(n421), .B(n408), .Z(n3405) );
  HS65_LL_NOR4ABX2 U12212 ( .A(n4672), .B(n4695), .C(n4543), .D(n4476), .Z(
        n4998) );
  HS65_LL_NOR4ABX2 U12213 ( .A(n6265), .B(n6288), .C(n6136), .D(n6069), .Z(
        n6591) );
  HS65_LL_NOR4ABX2 U12214 ( .A(n4833), .B(n4811), .C(n4620), .D(n4532), .Z(
        n5120) );
  HS65_LL_NOR4ABX2 U12215 ( .A(n6426), .B(n6404), .C(n6213), .D(n6125), .Z(
        n6712) );
  HS65_LL_CBI4I6X5 U12216 ( .A(n765), .B(n2052), .C(n785), .D(n2147), .Z(n2127) );
  HS65_LL_OA12X9 U12217 ( .A(n1970), .B(n790), .C(n769), .Z(n2147) );
  HS65_LL_CBI4I6X5 U12218 ( .A(n806), .B(n1676), .C(n826), .D(n1771), .Z(n1751) );
  HS65_LL_OA12X9 U12219 ( .A(n1594), .B(n831), .C(n810), .Z(n1771) );
  HS65_LL_NAND2X7 U12220 ( .A(n158), .B(n174), .Z(n3633) );
  HS65_LL_NAND2X7 U12221 ( .A(n17), .B(n31), .Z(n5105) );
  HS65_LL_NAND2X7 U12222 ( .A(n539), .B(n553), .Z(n6698) );
  HS65_LL_NAND4ABX3 U12223 ( .A(n6266), .B(n6267), .C(n6268), .D(n6269), .Z(
        n6066) );
  HS65_LL_NOR3AX2 U12224 ( .A(n6270), .B(n6271), .C(n6272), .Z(n6269) );
  HS65_LL_NAND3AX6 U12225 ( .A(n6273), .B(n6274), .C(n6275), .Z(n6267) );
  HS65_LL_AOI222X2 U12226 ( .A(n536), .B(n558), .C(n561), .D(n537), .E(n566), 
        .F(n538), .Z(n6268) );
  HS65_LL_NAND4ABX3 U12227 ( .A(n4673), .B(n4674), .C(n4675), .D(n4676), .Z(
        n4473) );
  HS65_LL_NOR3AX2 U12228 ( .A(n4677), .B(n4678), .C(n4679), .Z(n4676) );
  HS65_LL_NAND3AX6 U12229 ( .A(n4680), .B(n4681), .C(n4682), .Z(n4674) );
  HS65_LL_AOI222X2 U12230 ( .A(n14), .B(n36), .C(n39), .D(n15), .E(n44), .F(
        n16), .Z(n4675) );
  HS65_LL_NOR3AX2 U12231 ( .A(n4474), .B(n4543), .C(n4544), .Z(n4539) );
  HS65_LL_NOR3AX2 U12232 ( .A(n6067), .B(n6136), .C(n6137), .Z(n6132) );
  HS65_LL_NOR3AX2 U12233 ( .A(n4600), .B(n4767), .C(n4768), .Z(n4763) );
  HS65_LL_NOR3AX2 U12234 ( .A(n6193), .B(n6360), .C(n6361), .Z(n6356) );
  HS65_LL_NOR3AX2 U12235 ( .A(n6176), .B(n6321), .C(n6322), .Z(n6317) );
  HS65_LL_NOR3AX2 U12236 ( .A(n6123), .B(n6213), .C(n6214), .Z(n6209) );
  HS65_LL_NOR3AX2 U12237 ( .A(n4530), .B(n4620), .C(n4621), .Z(n4616) );
  HS65_LL_NAND2X7 U12238 ( .A(n157), .B(n173), .Z(n3255) );
  HS65_LL_NOR4ABX2 U12239 ( .A(n2986), .B(n2987), .C(n2988), .D(n2989), .Z(
        n2985) );
  HS65_LL_AO212X4 U12240 ( .A(n418), .B(n441), .C(n422), .D(n432), .E(n2990), 
        .Z(n2988) );
  HS65_LL_NAND2X7 U12241 ( .A(n60), .B(n74), .Z(n6488) );
  HS65_LL_NAND2X7 U12242 ( .A(n238), .B(n256), .Z(n4895) );
  HS65_LL_NAND2X7 U12243 ( .A(n499), .B(n510), .Z(n6413) );
  HS65_LL_NAND2X7 U12244 ( .A(n675), .B(n686), .Z(n4820) );
  HS65_LL_NOR2X6 U12245 ( .A(n122), .B(n134), .Z(n8832) );
  HS65_LL_NOR2X6 U12246 ( .A(n145), .B(n157), .Z(n3279) );
  HS65_LL_NOR3AX2 U12247 ( .A(n2906), .B(n3227), .C(n3020), .Z(n3221) );
  HS65_LL_NAND2X7 U12248 ( .A(n39), .B(n18), .Z(n5058) );
  HS65_LL_NAND2X7 U12249 ( .A(n561), .B(n540), .Z(n6651) );
  HS65_LL_NOR4ABX2 U12250 ( .A(n3647), .B(n3595), .C(n3608), .D(n3637), .Z(
        n4092) );
  HS65_LL_NOR3AX2 U12251 ( .A(n8069), .B(n7975), .C(n7856), .Z(n8064) );
  HS65_LL_NOR3AX2 U12252 ( .A(n7936), .B(n8043), .C(n8315), .Z(n8310) );
  HS65_LL_NOR2X6 U12253 ( .A(n319), .B(n325), .Z(n7770) );
  HS65_LL_NAND3X5 U12254 ( .A(n8810), .B(n8811), .C(n8812), .Z(n8439) );
  HS65_LL_NOR4ABX2 U12255 ( .A(n8817), .B(n7726), .C(n8818), .D(n7892), .Z(
        n8811) );
  HS65_LL_NOR4ABX2 U12256 ( .A(n8819), .B(n7925), .C(n8820), .D(n8821), .Z(
        n8810) );
  HS65_LL_NOR4ABX2 U12257 ( .A(n7912), .B(n8813), .C(n8814), .D(n8815), .Z(
        n8812) );
  HS65_LL_NOR2X6 U12258 ( .A(n365), .B(n374), .Z(n7752) );
  HS65_LL_NAND2X7 U12259 ( .A(n542), .B(n553), .Z(n6274) );
  HS65_LL_NAND2X7 U12260 ( .A(n20), .B(n31), .Z(n4681) );
  HS65_LL_NAND2X7 U12261 ( .A(n430), .B(n419), .Z(n3816) );
  HS65_LL_NOR2X6 U12262 ( .A(n47), .B(n33), .Z(n5113) );
  HS65_LL_NOR2X6 U12263 ( .A(n569), .B(n555), .Z(n6706) );
  HS65_LL_CBI4I6X5 U12264 ( .A(n475), .B(n477), .C(n455), .D(n5441), .Z(n5635)
         );
  HS65_LL_CBI4I6X5 U12265 ( .A(n684), .B(n690), .C(n675), .D(n5210), .Z(n5580)
         );
  HS65_LL_CBI4I6X5 U12266 ( .A(n508), .B(n514), .C(n499), .D(n6802), .Z(n7172)
         );
  HS65_LL_CBI4I6X5 U12267 ( .A(n300), .B(n302), .C(n280), .D(n7033), .Z(n7227)
         );
  HS65_LL_CBI4I6X5 U12268 ( .A(n258), .B(n260), .C(n238), .D(n5326), .Z(n5609)
         );
  HS65_LL_CBI4I6X5 U12269 ( .A(n73), .B(n83), .C(n60), .D(n6918), .Z(n7201) );
  HS65_LL_NAND2X7 U12270 ( .A(n120), .B(n106), .Z(n7909) );
  HS65_LL_NAND2X7 U12271 ( .A(n600), .B(n586), .Z(n7811) );
  HS65_LL_CBI4I6X5 U12272 ( .A(n29), .B(n35), .C(n20), .D(n5104), .Z(n5515) );
  HS65_LL_CBI4I6X5 U12273 ( .A(n551), .B(n557), .C(n542), .D(n6697), .Z(n7107)
         );
  HS65_LL_NOR2X6 U12274 ( .A(n469), .B(n474), .Z(n5449) );
  HS65_LL_NOR2X6 U12275 ( .A(n702), .B(n688), .Z(n5219) );
  HS65_LL_NOR2X6 U12276 ( .A(n526), .B(n512), .Z(n6811) );
  HS65_LL_NOR2X6 U12277 ( .A(n294), .B(n299), .Z(n7041) );
  HS65_LL_NOR2X6 U12278 ( .A(n252), .B(n257), .Z(n5334) );
  HS65_LL_NOR2X6 U12279 ( .A(n89), .B(n76), .Z(n6926) );
  HS65_LL_NOR2X6 U12280 ( .A(n180), .B(n166), .Z(n3575) );
  HS65_LL_NAND2X7 U12281 ( .A(n211), .B(n191), .Z(n3459) );
  HS65_LL_NOR2X6 U12282 ( .A(n344), .B(n355), .Z(n8528) );
  HS65_LL_NAND2X7 U12283 ( .A(n375), .B(n383), .Z(n8199) );
  HS65_LL_NOR2X6 U12284 ( .A(n812), .B(n803), .Z(n1744) );
  HS65_LL_NOR3AX2 U12285 ( .A(n6426), .B(n6121), .C(n6427), .Z(n6420) );
  HS65_LL_NOR3AX2 U12286 ( .A(n4833), .B(n4528), .C(n4834), .Z(n4827) );
  HS65_LL_NOR3AX2 U12287 ( .A(n8325), .B(n7939), .C(n8326), .Z(n8318) );
  HS65_LL_NOR3AX2 U12288 ( .A(n6404), .B(n6214), .C(n6122), .Z(n6399) );
  HS65_LL_NOR3AX2 U12289 ( .A(n4811), .B(n4621), .C(n4529), .Z(n4806) );
  HS65_LL_NOR3AX2 U12290 ( .A(n3170), .B(n3171), .C(n2989), .Z(n3166) );
  HS65_LL_NOR2X6 U12291 ( .A(n226), .B(n221), .Z(n3451) );
  HS65_LL_NOR2X6 U12292 ( .A(n383), .B(n393), .Z(n8303) );
  HS65_LL_NOR4ABX2 U12293 ( .A(n8220), .B(n8221), .C(n8222), .D(n8223), .Z(
        n8214) );
  HS65_LL_NAND2X7 U12294 ( .A(n629), .B(n645), .Z(n3664) );
  HS65_LL_NOR2X6 U12295 ( .A(n645), .B(n650), .Z(n3693) );
  HS65_LL_NOR3AX2 U12296 ( .A(n8376), .B(n7999), .C(n8140), .Z(n8372) );
  HS65_LL_NOR3AX2 U12297 ( .A(n8428), .B(n8012), .C(n8163), .Z(n8424) );
  HS65_LL_NOR2X6 U12298 ( .A(n432), .B(n441), .Z(n3808) );
  HS65_LL_NAND2X7 U12299 ( .A(n197), .B(n226), .Z(n3421) );
  HS65_LL_NAND2X7 U12300 ( .A(n152), .B(n180), .Z(n3545) );
  HS65_LL_NOR3AX2 U12301 ( .A(n3495), .B(n2951), .C(n3531), .Z(n4065) );
  HS65_LL_NAND2X7 U12302 ( .A(n590), .B(n603), .Z(n8676) );
  HS65_LL_NAND2X7 U12303 ( .A(n143), .B(n177), .Z(n2920) );
  HS65_LL_NOR4ABX2 U12304 ( .A(n8392), .B(n7687), .C(n7799), .D(n8393), .Z(
        n8391) );
  HS65_LL_NOR4ABX2 U12305 ( .A(n8444), .B(n7725), .C(n7898), .D(n8445), .Z(
        n8443) );
  HS65_LL_NOR4ABX2 U12306 ( .A(n3482), .B(n3483), .C(n3484), .D(n3485), .Z(
        n3481) );
  HS65_LL_NOR4ABX2 U12307 ( .A(n6812), .B(n6813), .C(n6814), .D(n6815), .Z(
        n6426) );
  HS65_LL_NAND3AX6 U12308 ( .A(n6816), .B(n6817), .C(n6818), .Z(n6814) );
  HS65_LL_MX41X7 U12309 ( .D0(n494), .S0(n520), .D1(n524), .S1(n498), .D2(n508), .S2(n496), .D3(n513), .S3(n497), .Z(n6815) );
  HS65_LL_NOR4ABX2 U12310 ( .A(n6824), .B(n6825), .C(n6826), .D(n6827), .Z(
        n6812) );
  HS65_LL_NOR4ABX2 U12311 ( .A(n5220), .B(n5221), .C(n5222), .D(n5223), .Z(
        n4833) );
  HS65_LL_NAND3AX6 U12312 ( .A(n5224), .B(n5225), .C(n5226), .Z(n5222) );
  HS65_LL_MX41X7 U12313 ( .D0(n670), .S0(n696), .D1(n700), .S1(n674), .D2(n684), .S2(n672), .D3(n689), .S3(n673), .Z(n5223) );
  HS65_LL_NOR4ABX2 U12314 ( .A(n5232), .B(n5233), .C(n5234), .D(n5235), .Z(
        n5220) );
  HS65_LL_NOR4ABX2 U12315 ( .A(n5100), .B(n5101), .C(n5102), .D(n5103), .Z(
        n4672) );
  HS65_LL_NAND3AX6 U12316 ( .A(n5104), .B(n5105), .C(n5106), .Z(n5103) );
  HS65_LL_NAND4ABX3 U12317 ( .A(n5107), .B(n5108), .C(n5109), .D(n5110), .Z(
        n5102) );
  HS65_LL_AOI222X2 U12318 ( .A(n39), .B(n9), .C(n33), .D(n4569), .E(n10), .F(
        n30), .Z(n5100) );
  HS65_LL_NOR4ABX2 U12319 ( .A(n6693), .B(n6694), .C(n6695), .D(n6696), .Z(
        n6265) );
  HS65_LL_NAND3AX6 U12320 ( .A(n6697), .B(n6698), .C(n6699), .Z(n6696) );
  HS65_LL_NAND4ABX3 U12321 ( .A(n6700), .B(n6701), .C(n6702), .D(n6703), .Z(
        n6695) );
  HS65_LL_AOI222X2 U12322 ( .A(n561), .B(n531), .C(n555), .D(n6162), .E(n532), 
        .F(n552), .Z(n6693) );
  HS65_LL_NOR4ABX2 U12323 ( .A(n8595), .B(n8596), .C(n8597), .D(n8598), .Z(
        n8325) );
  HS65_LL_NAND4ABX3 U12324 ( .A(n8599), .B(n8600), .C(n8601), .D(n8602), .Z(
        n8597) );
  HS65_LL_MX41X7 U12325 ( .D0(n332), .S0(n340), .D1(n323), .S1(n345), .D2(n353), .S2(n334), .D3(n324), .S3(n349), .Z(n8598) );
  HS65_LL_NOR3AX2 U12326 ( .A(n8603), .B(n8604), .C(n8605), .Z(n8596) );
  HS65_LL_NAND2X7 U12327 ( .A(n340), .B(n326), .Z(n8578) );
  HS65_LL_NOR3AX2 U12328 ( .A(n3850), .B(n3178), .C(n3885), .Z(n4312) );
  HS65_LL_NOR3AX2 U12329 ( .A(n3735), .B(n3152), .C(n3770), .Z(n4253) );
  HS65_LL_NOR4ABX2 U12330 ( .A(n8102), .B(n8103), .C(n8104), .D(n8105), .Z(
        n8096) );
  HS65_LL_NAND2X7 U12331 ( .A(n152), .B(n165), .Z(n3038) );
  HS65_LL_NOR4ABX2 U12332 ( .A(n3652), .B(n3606), .C(n3594), .D(n3631), .Z(
        n4122) );
  HS65_LL_NAND2X7 U12333 ( .A(n612), .B(n593), .Z(n8751) );
  HS65_LL_NAND2X7 U12334 ( .A(n18), .B(n35), .Z(n5032) );
  HS65_LL_NAND2X7 U12335 ( .A(n540), .B(n557), .Z(n6625) );
  HS65_LL_NOR4ABX2 U12336 ( .A(n5322), .B(n5323), .C(n5324), .D(n5325), .Z(
        n4886) );
  HS65_LL_NAND3AX6 U12337 ( .A(n5326), .B(n5327), .C(n5328), .Z(n5325) );
  HS65_LL_NAND4ABX3 U12338 ( .A(n5329), .B(n5330), .C(n5331), .D(n5332), .Z(
        n5324) );
  HS65_LL_AOI222X2 U12339 ( .A(n245), .B(n268), .C(n257), .D(n4730), .E(n247), 
        .F(n259), .Z(n5322) );
  HS65_LL_NOR4ABX2 U12340 ( .A(n5437), .B(n5438), .C(n5439), .D(n5440), .Z(
        n4939) );
  HS65_LL_NAND3AX6 U12341 ( .A(n5441), .B(n5442), .C(n5443), .Z(n5440) );
  HS65_LL_NAND4ABX3 U12342 ( .A(n5444), .B(n5445), .C(n5446), .D(n5447), .Z(
        n5439) );
  HS65_LL_AOI222X2 U12343 ( .A(n462), .B(n485), .C(n474), .D(n4792), .E(n464), 
        .F(n476), .Z(n5437) );
  HS65_LL_NOR4ABX2 U12344 ( .A(n5206), .B(n5207), .C(n5208), .D(n5209), .Z(
        n4811) );
  HS65_LL_NAND3AX6 U12345 ( .A(n5210), .B(n5211), .C(n5212), .Z(n5209) );
  HS65_LL_NAND4ABX3 U12346 ( .A(n5213), .B(n5214), .C(n5215), .D(n5216), .Z(
        n5208) );
  HS65_LL_AOI222X2 U12347 ( .A(n665), .B(n694), .C(n688), .D(n4646), .E(n666), 
        .F(n685), .Z(n5206) );
  HS65_LL_NOR4ABX2 U12348 ( .A(n7029), .B(n7030), .C(n7031), .D(n7032), .Z(
        n6532) );
  HS65_LL_NAND3AX6 U12349 ( .A(n7033), .B(n7034), .C(n7035), .Z(n7032) );
  HS65_LL_NAND4ABX3 U12350 ( .A(n7036), .B(n7037), .C(n7038), .D(n7039), .Z(
        n7031) );
  HS65_LL_AOI222X2 U12351 ( .A(n287), .B(n310), .C(n299), .D(n6385), .E(n289), 
        .F(n301), .Z(n7029) );
  HS65_LL_NOR4ABX2 U12352 ( .A(n6798), .B(n6799), .C(n6800), .D(n6801), .Z(
        n6404) );
  HS65_LL_NAND3AX6 U12353 ( .A(n6802), .B(n6803), .C(n6804), .Z(n6801) );
  HS65_LL_NAND4ABX3 U12354 ( .A(n6805), .B(n6806), .C(n6807), .D(n6808), .Z(
        n6800) );
  HS65_LL_AOI222X2 U12355 ( .A(n489), .B(n518), .C(n512), .D(n6239), .E(n490), 
        .F(n509), .Z(n6798) );
  HS65_LL_NOR4ABX2 U12356 ( .A(n6755), .B(n6756), .C(n6757), .D(n6758), .Z(
        n6749) );
  HS65_LL_NOR4ABX2 U12357 ( .A(n5163), .B(n5164), .C(n5165), .D(n5166), .Z(
        n5157) );
  HS65_LL_NOR4ABX2 U12358 ( .A(n5395), .B(n5396), .C(n5397), .D(n5398), .Z(
        n5389) );
  HS65_LL_NAND2X7 U12359 ( .A(n673), .B(n690), .Z(n5154) );
  HS65_LL_NAND2X7 U12360 ( .A(n497), .B(n514), .Z(n6746) );
  HS65_LL_NAND2X7 U12361 ( .A(n197), .B(n224), .Z(n3420) );
  HS65_LL_NOR4ABX2 U12362 ( .A(n8822), .B(n8823), .C(n8824), .D(n8825), .Z(
        n8428) );
  HS65_LL_NAND3AX6 U12363 ( .A(n8826), .B(n7906), .C(n8827), .Z(n8825) );
  HS65_LL_NAND4ABX3 U12364 ( .A(n8828), .B(n8829), .C(n8830), .D(n7893), .Z(
        n8824) );
  HS65_LL_AOI222X2 U12365 ( .A(n104), .B(n129), .C(n134), .D(n8181), .E(n103), 
        .F(n136), .Z(n8822) );
  HS65_LL_NOR4ABX2 U12366 ( .A(n3875), .B(n3831), .C(n3847), .D(n3866), .Z(
        n4300) );
  HS65_LL_NOR4ABX2 U12367 ( .A(n3247), .B(n3248), .C(n3249), .D(n3250), .Z(
        n3241) );
  HS65_LL_NOR4ABX2 U12368 ( .A(n4971), .B(n4972), .C(n4973), .D(n4974), .Z(
        n4965) );
  HS65_LL_NOR4ABX2 U12369 ( .A(n6436), .B(n6437), .C(n6438), .D(n6439), .Z(
        n6430) );
  HS65_LL_NOR4ABX2 U12370 ( .A(n4843), .B(n4844), .C(n4845), .D(n4846), .Z(
        n4837) );
  HS65_LL_NOR4ABX2 U12371 ( .A(n3453), .B(n3454), .C(n3455), .D(n3456), .Z(
        n2943) );
  HS65_LL_NAND4ABX3 U12372 ( .A(n3457), .B(n3458), .C(n3459), .D(n3460), .Z(
        n3456) );
  HS65_LL_AOI212X4 U12373 ( .A(n224), .B(n3461), .C(n213), .D(n3462), .E(n3463), .Z(n3454) );
  HS65_LL_MX41X7 U12374 ( .D0(n198), .S0(n226), .D1(n219), .S1(n203), .D2(n215), .S2(n191), .D3(n211), .S3(n196), .Z(n3455) );
  HS65_LL_NOR4ABX2 U12375 ( .A(n3577), .B(n3578), .C(n3579), .D(n3580), .Z(
        n3019) );
  HS65_LL_NAND4ABX3 U12376 ( .A(n3581), .B(n3582), .C(n3583), .D(n3584), .Z(
        n3580) );
  HS65_LL_MX41X7 U12377 ( .D0(n153), .S0(n180), .D1(n158), .S1(n164), .D2(n170), .S2(n146), .D3(n175), .S3(n151), .Z(n3579) );
  HS65_LL_AOI212X4 U12378 ( .A(n178), .B(n3585), .C(n167), .D(n3586), .E(n3587), .Z(n3578) );
  HS65_LL_NOR4ABX2 U12379 ( .A(n8335), .B(n8336), .C(n8337), .D(n8338), .Z(
        n8329) );
  HS65_LL_NOR4ABX2 U12380 ( .A(n3810), .B(n3811), .C(n3812), .D(n3813), .Z(
        n3170) );
  HS65_LL_NAND4ABX3 U12381 ( .A(n3814), .B(n3815), .C(n3816), .D(n3817), .Z(
        n3813) );
  HS65_LL_MX41X7 U12382 ( .D0(n413), .S0(n432), .D1(n442), .S1(n406), .D2(n437), .S2(n419), .D3(n430), .S3(n409), .Z(n3812) );
  HS65_LL_AOI212X4 U12383 ( .A(n433), .B(n3818), .C(n439), .D(n3819), .E(n3820), .Z(n3811) );
  HS65_LL_NOR4ABX2 U12384 ( .A(n3695), .B(n3696), .C(n3697), .D(n3698), .Z(
        n3144) );
  HS65_LL_NAND4ABX3 U12385 ( .A(n3699), .B(n3700), .C(n3701), .D(n3702), .Z(
        n3698) );
  HS65_LL_MX41X7 U12386 ( .D0(n631), .S0(n645), .D1(n651), .S1(n625), .D2(n654), .S2(n637), .D3(n661), .S3(n628), .Z(n3697) );
  HS65_LL_AOI222X2 U12387 ( .A(n633), .B(n658), .C(n626), .D(n649), .E(n636), 
        .F(n660), .Z(n3695) );
  HS65_LL_NOR3AX2 U12388 ( .A(n3685), .B(n3686), .C(n3687), .Z(n3684) );
  HS65_LL_NAND4ABX3 U12389 ( .A(n8543), .B(n8544), .C(n8545), .D(n8546), .Z(
        n8041) );
  HS65_LL_NOR3AX2 U12390 ( .A(n8551), .B(n8552), .C(n8553), .Z(n8545) );
  HS65_LL_NAND4ABX3 U12391 ( .A(n8557), .B(n8558), .C(n7762), .D(n8559), .Z(
        n8543) );
  HS65_LL_NOR4ABX2 U12392 ( .A(n8547), .B(n8548), .C(n8549), .D(n8550), .Z(
        n8546) );
  HS65_LL_NAND4ABX3 U12393 ( .A(n3602), .B(n3603), .C(n3604), .D(n3605), .Z(
        n3018) );
  HS65_LL_NOR3AX2 U12394 ( .A(n3610), .B(n3611), .C(n3612), .Z(n3604) );
  HS65_LL_NOR4ABX2 U12395 ( .A(n3606), .B(n3607), .C(n3608), .D(n3609), .Z(
        n3605) );
  HS65_LL_NAND4ABX3 U12396 ( .A(n3616), .B(n3617), .C(n3618), .D(n3619), .Z(
        n3602) );
  HS65_LL_NAND4ABX3 U12397 ( .A(n6607), .B(n6608), .C(n6609), .D(n6610), .Z(
        n6135) );
  HS65_LL_NOR3X4 U12398 ( .A(n6615), .B(n6616), .C(n6617), .Z(n6609) );
  HS65_LL_NOR4ABX2 U12399 ( .A(n6611), .B(n6612), .C(n6613), .D(n6614), .Z(
        n6610) );
  HS65_LL_NAND4ABX3 U12400 ( .A(n6622), .B(n6623), .C(n6624), .D(n6625), .Z(
        n6607) );
  HS65_LL_NAND4ABX3 U12401 ( .A(n5014), .B(n5015), .C(n5016), .D(n5017), .Z(
        n4542) );
  HS65_LL_NOR3X4 U12402 ( .A(n5022), .B(n5023), .C(n5024), .Z(n5016) );
  HS65_LL_NOR4ABX2 U12403 ( .A(n5018), .B(n5019), .C(n5020), .D(n5021), .Z(
        n5017) );
  HS65_LL_NAND4ABX3 U12404 ( .A(n5029), .B(n5030), .C(n5031), .D(n5032), .Z(
        n5014) );
  HS65_LL_NAND2X7 U12405 ( .A(n398), .B(n365), .Z(n7986) );
  HS65_LL_NAND2X7 U12406 ( .A(n459), .B(n469), .Z(n5385) );
  HS65_LL_NAND2X7 U12407 ( .A(n242), .B(n252), .Z(n5270) );
  HS65_LL_NAND2X7 U12408 ( .A(n284), .B(n294), .Z(n6977) );
  HS65_LL_NAND2X7 U12409 ( .A(n671), .B(n702), .Z(n5153) );
  HS65_LL_NAND2X7 U12410 ( .A(n495), .B(n526), .Z(n6745) );
  HS65_LL_NAND2X7 U12411 ( .A(n152), .B(n169), .Z(n3576) );
  HS65_LL_NAND2X7 U12412 ( .A(n462), .B(n474), .Z(n5404) );
  HS65_LL_NAND2X7 U12413 ( .A(n287), .B(n299), .Z(n6996) );
  HS65_LL_NAND2X7 U12414 ( .A(n665), .B(n688), .Z(n5173) );
  HS65_LL_NAND2X7 U12415 ( .A(n489), .B(n512), .Z(n6765) );
  HS65_LL_NAND2X7 U12416 ( .A(n191), .B(n226), .Z(n3515) );
  HS65_LL_NAND4ABX3 U12417 ( .A(n4089), .B(n4090), .C(n4091), .D(n4092), .Z(
        n3906) );
  HS65_LL_AOI222X2 U12418 ( .A(n142), .B(n163), .C(n152), .D(n170), .E(n164), 
        .F(n157), .Z(n4091) );
  HS65_LL_NAND4ABX3 U12419 ( .A(n3569), .B(n3553), .C(n4094), .D(n3584), .Z(
        n4089) );
  HS65_LL_NAND4ABX3 U12420 ( .A(n3276), .B(n3260), .C(n3026), .D(n3244), .Z(
        n4090) );
  HS65_LL_OAI21X3 U12421 ( .A(n285), .B(n6543), .C(n292), .Z(n6542) );
  HS65_LL_OAI21X3 U12422 ( .A(n56), .B(n6490), .C(n91), .Z(n6489) );
  HS65_LL_OAI21X3 U12423 ( .A(n243), .B(n4897), .C(n250), .Z(n4896) );
  HS65_LL_OAI21X3 U12424 ( .A(n460), .B(n4950), .C(n467), .Z(n4949) );
  HS65_LL_OAI21X3 U12425 ( .A(n496), .B(n6415), .C(n525), .Z(n6414) );
  HS65_LL_OAI21X3 U12426 ( .A(n672), .B(n4822), .C(n701), .Z(n4821) );
  HS65_LL_NAND2X7 U12427 ( .A(n106), .B(n122), .Z(n8758) );
  HS65_LL_NAND2X7 U12428 ( .A(n586), .B(n602), .Z(n8668) );
  HS65_LL_OAI21X3 U12429 ( .A(n450), .B(n4950), .C(n484), .Z(n5560) );
  HS65_LL_OAI21X3 U12430 ( .A(n233), .B(n4897), .C(n267), .Z(n5538) );
  HS65_LL_OAI21X3 U12431 ( .A(n678), .B(n4822), .C(n696), .Z(n5495) );
  HS65_LL_OAI21X3 U12432 ( .A(n275), .B(n6543), .C(n309), .Z(n7152) );
  HS65_LL_OAI21X3 U12433 ( .A(n502), .B(n6415), .C(n520), .Z(n7087) );
  HS65_LL_OAI21X3 U12434 ( .A(n64), .B(n6490), .C(n81), .Z(n7130) );
  HS65_LL_NAND2X7 U12435 ( .A(n64), .B(n89), .Z(n6834) );
  HS65_LL_NAND2X7 U12436 ( .A(n233), .B(n252), .Z(n5242) );
  HS65_LL_NAND2X7 U12437 ( .A(n450), .B(n469), .Z(n5357) );
  HS65_LL_NAND2X7 U12438 ( .A(n678), .B(n702), .Z(n5124) );
  HS65_LL_NAND2X7 U12439 ( .A(n275), .B(n294), .Z(n6949) );
  HS65_LL_NAND2X7 U12440 ( .A(n502), .B(n526), .Z(n6716) );
  HS65_LL_NAND2X7 U12441 ( .A(n23), .B(n35), .Z(n5110) );
  HS65_LL_NAND2X7 U12442 ( .A(n545), .B(n557), .Z(n6703) );
  HS65_LL_NAND2X7 U12443 ( .A(n146), .B(n178), .Z(n3244) );
  HS65_LL_NAND2X7 U12444 ( .A(n391), .B(n375), .Z(n8122) );
  HS65_LL_NAND2X7 U12445 ( .A(n327), .B(n344), .Z(n8502) );
  HS65_LL_NAND2X7 U12446 ( .A(n329), .B(n355), .Z(n7762) );
  HS65_LL_NAND2X7 U12447 ( .A(n108), .B(n125), .Z(n7907) );
  HS65_LL_NAND2X7 U12448 ( .A(n588), .B(n605), .Z(n7809) );
  HS65_LL_OAI21X3 U12449 ( .A(n370), .B(n8080), .C(n387), .Z(n8079) );
  HS65_LL_OAI21X3 U12450 ( .A(n334), .B(n8324), .C(n348), .Z(n8355) );
  HS65_LL_NAND2X7 U12451 ( .A(n64), .B(n83), .Z(n6923) );
  HS65_LL_NAND2X7 U12452 ( .A(n233), .B(n260), .Z(n5331) );
  HS65_LL_NAND2X7 U12453 ( .A(n450), .B(n477), .Z(n5446) );
  HS65_LL_NAND2X7 U12454 ( .A(n678), .B(n690), .Z(n5215) );
  HS65_LL_NAND2X7 U12455 ( .A(n275), .B(n302), .Z(n7038) );
  HS65_LL_NAND2X7 U12456 ( .A(n502), .B(n514), .Z(n6807) );
  HS65_LL_NAND2X7 U12457 ( .A(n166), .B(n157), .Z(n3647) );
  HS65_LL_NAND2X7 U12458 ( .A(n604), .B(n582), .Z(n8148) );
  HS65_LL_NAND2X7 U12459 ( .A(n124), .B(n102), .Z(n8171) );
  HS65_LL_OAI21X3 U12460 ( .A(n629), .B(n3311), .C(n659), .Z(n3936) );
  HS65_LL_OAI21X3 U12461 ( .A(n375), .B(n8080), .C(n389), .Z(n8482) );
  HS65_LL_NAND2X7 U12462 ( .A(n329), .B(n351), .Z(n8529) );
  HS65_LL_OAI21X3 U12463 ( .A(n327), .B(n8324), .C(n340), .Z(n8872) );
  HS65_LL_NAND2X7 U12464 ( .A(n23), .B(n47), .Z(n5003) );
  HS65_LL_NAND2X7 U12465 ( .A(n545), .B(n569), .Z(n6596) );
  HS65_LL_NOR2X6 U12466 ( .A(n288), .B(n282), .Z(n6580) );
  HS65_LL_NOR2X6 U12467 ( .A(n67), .B(n62), .Z(n6468) );
  HS65_LL_NOR2X6 U12468 ( .A(n246), .B(n240), .Z(n4875) );
  HS65_LL_NOR2X6 U12469 ( .A(n463), .B(n457), .Z(n4987) );
  HS65_LL_NOR2X6 U12470 ( .A(n492), .B(n500), .Z(n6454) );
  HS65_LL_NOR2X6 U12471 ( .A(n668), .B(n676), .Z(n4861) );
  HS65_LL_NAND2X7 U12472 ( .A(n147), .B(n169), .Z(n3551) );
  HS65_LL_NAND2X7 U12473 ( .A(n197), .B(n211), .Z(n3430) );
  HS65_LL_NOR2X6 U12474 ( .A(n582), .B(n590), .Z(n7677) );
  HS65_LL_NOR2X6 U12475 ( .A(n102), .B(n110), .Z(n7715) );
  HS65_LL_OAI21X3 U12476 ( .A(n586), .B(n8385), .C(n610), .Z(n9052) );
  HS65_LL_OAI21X3 U12477 ( .A(n106), .B(n8437), .C(n130), .Z(n9110) );
  HS65_LL_NAND2X7 U12478 ( .A(n437), .B(n415), .Z(n3388) );
  HS65_LL_NAND2X7 U12479 ( .A(n215), .B(n192), .Z(n3105) );
  HS65_LL_NAND2X7 U12480 ( .A(n579), .B(n610), .Z(n7790) );
  HS65_LL_NAND2X7 U12481 ( .A(n99), .B(n130), .Z(n7889) );
  HS65_LL_NAND2X7 U12482 ( .A(n524), .B(n497), .Z(n6786) );
  HS65_LL_NAND2X7 U12483 ( .A(n700), .B(n673), .Z(n5194) );
  HS65_LL_NAND2X7 U12484 ( .A(n23), .B(n42), .Z(n5093) );
  HS65_LL_NAND2X7 U12485 ( .A(n545), .B(n564), .Z(n6686) );
  HS65_LL_NAND2X7 U12486 ( .A(n197), .B(n210), .Z(n3066) );
  HS65_LL_NAND2X7 U12487 ( .A(n411), .B(n429), .Z(n3411) );
  HS65_LL_NAND2X7 U12488 ( .A(n108), .B(n137), .Z(n7908) );
  HS65_LL_NAND2X7 U12489 ( .A(n588), .B(n617), .Z(n7810) );
  HS65_LL_NAND2X7 U12490 ( .A(n363), .B(n391), .Z(n8107) );
  HS65_LL_OAI21X3 U12491 ( .A(n865), .B(n868), .C(n854), .Z(n1122) );
  HS65_LL_OAI21X3 U12492 ( .A(n783), .B(n786), .C(n772), .Z(n1874) );
  HS65_LL_OAI21X3 U12493 ( .A(n14), .B(n9), .C(n30), .Z(n5756) );
  HS65_LL_OAI21X3 U12494 ( .A(n536), .B(n531), .C(n552), .Z(n7348) );
  HS65_LL_OAI21X3 U12495 ( .A(n539), .B(n6276), .C(n568), .Z(n6275) );
  HS65_LL_OAI21X3 U12496 ( .A(n17), .B(n4683), .C(n46), .Z(n4682) );
  HS65_LL_NAND2X7 U12497 ( .A(n147), .B(n174), .Z(n3025) );
  HS65_LL_IVX9 U12498 ( .A(n2795), .Z(n230) );
  HS65_LL_OAI21X3 U12499 ( .A(n824), .B(n827), .C(n813), .Z(n1498) );
  HS65_LL_NAND2X7 U12500 ( .A(n192), .B(n220), .Z(n3494) );
  HS65_LL_NAND2X7 U12501 ( .A(n112), .B(n131), .Z(n7708) );
  HS65_LL_NAND2X7 U12502 ( .A(n174), .B(n157), .Z(n3646) );
  HS65_LL_OAI21X3 U12503 ( .A(n906), .B(n909), .C(n895), .Z(n2250) );
  HS65_LL_NAND2X7 U12504 ( .A(n126), .B(n108), .Z(n7893) );
  HS65_LL_NAND2X7 U12505 ( .A(n606), .B(n588), .Z(n7794) );
  HS65_LL_NAND3AX6 U12506 ( .A(n3098), .B(n3099), .C(n3100), .Z(n3083) );
  HS65_LL_AOI12X2 U12507 ( .A(n188), .B(n3101), .C(n3102), .Z(n3100) );
  HS65_LL_NAND2X7 U12508 ( .A(n325), .B(n349), .Z(n8577) );
  HS65_LL_OAI21X3 U12509 ( .A(n672), .B(n669), .C(n699), .Z(n5766) );
  HS65_LL_OAI21X3 U12510 ( .A(n23), .B(n4683), .C(n41), .Z(n5471) );
  HS65_LL_OAI21X3 U12511 ( .A(n545), .B(n6276), .C(n563), .Z(n7063) );
  HS65_LL_OAI21X3 U12512 ( .A(n411), .B(n3365), .C(n428), .Z(n3974) );
  HS65_LL_OAI21X3 U12513 ( .A(n197), .B(n3080), .C(n212), .Z(n3891) );
  HS65_LL_NAND2X7 U12514 ( .A(n165), .B(n150), .Z(n3629) );
  HS65_LL_IVX9 U12515 ( .A(n2779), .Z(n572) );
  HS65_LL_OAI21X3 U12516 ( .A(n192), .B(n188), .C(n219), .Z(n4225) );
  HS65_LL_NAND2X7 U12517 ( .A(n152), .B(n173), .Z(n3285) );
  HS65_LL_NAND2X7 U12518 ( .A(n829), .B(n804), .Z(n1559) );
  HS65_LL_AOI12X2 U12519 ( .A(n552), .B(n541), .C(n6653), .Z(n6652) );
  HS65_LL_AOI12X2 U12520 ( .A(n30), .B(n19), .C(n5060), .Z(n5059) );
  HS65_LL_NAND2X7 U12521 ( .A(n367), .B(n400), .Z(n8226) );
  HS65_LL_OAI21X3 U12522 ( .A(n175), .B(n3040), .C(n156), .Z(n3039) );
  HS65_LL_NAND2X7 U12523 ( .A(n190), .B(n220), .Z(n3431) );
  HS65_LL_NAND2X7 U12524 ( .A(n421), .B(n440), .Z(n3789) );
  HS65_LL_NAND2X7 U12525 ( .A(n412), .B(n438), .Z(n3188) );
  HS65_LL_NAND2X7 U12526 ( .A(n586), .B(n611), .Z(n8420) );
  HS65_LL_NAND2X7 U12527 ( .A(n106), .B(n131), .Z(n8472) );
  HS65_LL_AOI12X2 U12528 ( .A(n170), .B(n150), .C(n3561), .Z(n3560) );
  HS65_LL_NAND2X7 U12529 ( .A(n633), .B(n653), .Z(n3678) );
  HS65_LL_NAND2X7 U12530 ( .A(n630), .B(n655), .Z(n3161) );
  HS65_LL_NAND2X7 U12531 ( .A(n422), .B(n429), .Z(n3382) );
  HS65_LL_NAND2X7 U12532 ( .A(n189), .B(n210), .Z(n3099) );
  HS65_LL_NAND2X7 U12533 ( .A(n178), .B(n155), .Z(n3595) );
  HS65_LL_NAND2X7 U12534 ( .A(n459), .B(n473), .Z(n5399) );
  HS65_LL_NAND2X7 U12535 ( .A(n284), .B(n298), .Z(n6991) );
  HS65_LL_NAND2X7 U12536 ( .A(n671), .B(n686), .Z(n5167) );
  HS65_LL_NAND2X7 U12537 ( .A(n495), .B(n510), .Z(n6759) );
  HS65_LL_OAI21X3 U12538 ( .A(n793), .B(n786), .C(n769), .Z(n1918) );
  HS65_LL_OAI21X3 U12539 ( .A(n10), .B(n9), .C(n41), .Z(n4575) );
  HS65_LL_OAI21X3 U12540 ( .A(n532), .B(n531), .C(n563), .Z(n6168) );
  HS65_LL_AOI12X2 U12541 ( .A(n478), .B(n459), .C(n5457), .Z(n5456) );
  HS65_LL_AOI12X2 U12542 ( .A(n516), .B(n495), .C(n6819), .Z(n6818) );
  HS65_LL_AOI12X2 U12543 ( .A(n692), .B(n671), .C(n5227), .Z(n5226) );
  HS65_LL_AOI12X2 U12544 ( .A(n322), .B(n8343), .C(n8344), .Z(n8342) );
  HS65_LL_NAND2X7 U12545 ( .A(n199), .B(n214), .Z(n2961) );
  HS65_LL_OAI21X3 U12546 ( .A(n834), .B(n827), .C(n810), .Z(n1542) );
  HS65_LL_NAND2X7 U12547 ( .A(n275), .B(n307), .Z(n6586) );
  HS65_LL_NAND2X7 U12548 ( .A(n233), .B(n265), .Z(n4881) );
  HS65_LL_NAND2X7 U12549 ( .A(n450), .B(n482), .Z(n4993) );
  HS65_LL_NAND2X7 U12550 ( .A(n502), .B(n519), .Z(n6460) );
  HS65_LL_NAND2X7 U12551 ( .A(n678), .B(n695), .Z(n4867) );
  HS65_LL_OAI21X3 U12552 ( .A(n916), .B(n909), .C(n892), .Z(n2294) );
  HS65_LL_AOI12X2 U12553 ( .A(n37), .B(n16), .C(n5091), .Z(n5090) );
  HS65_LL_AOI12X2 U12554 ( .A(n559), .B(n538), .C(n6684), .Z(n6683) );
  HS65_LL_NAND2X7 U12555 ( .A(n168), .B(n149), .Z(n3550) );
  HS65_LL_NAND2X7 U12556 ( .A(n154), .B(n173), .Z(n3571) );
  HS65_LL_NAND2X7 U12557 ( .A(n21), .B(n40), .Z(n4702) );
  HS65_LL_NAND2X7 U12558 ( .A(n543), .B(n562), .Z(n6295) );
  HS65_LL_NAND2X7 U12559 ( .A(n676), .B(n695), .Z(n4840) );
  HS65_LL_NAND2X7 U12560 ( .A(n500), .B(n519), .Z(n6433) );
  HS65_LL_NAND2X7 U12561 ( .A(n492), .B(n510), .Z(n6821) );
  HS65_LL_NAND2X7 U12562 ( .A(n668), .B(n686), .Z(n5229) );
  HS65_LL_OAI21X3 U12563 ( .A(n189), .B(n188), .C(n212), .Z(n2936) );
  HS65_LL_AOI12X2 U12564 ( .A(n509), .B(n498), .C(n6774), .Z(n6773) );
  HS65_LL_AOI12X2 U12565 ( .A(n685), .B(n674), .C(n5182), .Z(n5181) );
  HS65_LL_AOI12X2 U12566 ( .A(n476), .B(n453), .C(n5413), .Z(n5412) );
  HS65_LL_NAND2X7 U12567 ( .A(n16), .B(n31), .Z(n5045) );
  HS65_LL_NAND2X7 U12568 ( .A(n538), .B(n553), .Z(n6638) );
  HS65_LL_OAI21X3 U12569 ( .A(n37), .B(n29), .C(n18), .Z(n4666) );
  HS65_LL_OAI21X3 U12570 ( .A(n559), .B(n551), .C(n540), .Z(n6259) );
  HS65_LL_AOI12X2 U12571 ( .A(n566), .B(n546), .C(n6641), .Z(n6640) );
  HS65_LL_AOI12X2 U12572 ( .A(n44), .B(n24), .C(n5048), .Z(n5047) );
  HS65_LL_OAI21X3 U12573 ( .A(n390), .B(n397), .C(n368), .Z(n8994) );
  HS65_LL_NAND2X7 U12574 ( .A(n463), .B(n472), .Z(n5396) );
  HS65_LL_NAND2X7 U12575 ( .A(n288), .B(n297), .Z(n6988) );
  HS65_LL_NAND2X7 U12576 ( .A(n668), .B(n699), .Z(n5164) );
  HS65_LL_NAND2X7 U12577 ( .A(n492), .B(n523), .Z(n6756) );
  HS65_LL_OAI21X3 U12578 ( .A(n485), .B(n479), .C(n459), .Z(n5637) );
  HS65_LL_OAI21X3 U12579 ( .A(n310), .B(n304), .C(n284), .Z(n7229) );
  HS65_LL_OAI21X3 U12580 ( .A(n268), .B(n262), .C(n242), .Z(n5589) );
  HS65_LL_OAI21X3 U12581 ( .A(n82), .B(n84), .C(n54), .Z(n7181) );
  HS65_LL_OAI21X3 U12582 ( .A(n518), .B(n515), .C(n495), .Z(n7175) );
  HS65_LL_OAI21X3 U12583 ( .A(n694), .B(n691), .C(n671), .Z(n5583) );
  HS65_LL_OAI21X3 U12584 ( .A(n167), .B(n175), .C(n156), .Z(n4156) );
  HS65_LL_NAND2X7 U12585 ( .A(n329), .B(n347), .Z(n8564) );
  HS65_LL_OAI21X3 U12586 ( .A(n213), .B(n211), .C(n201), .Z(n4190) );
  HS65_LL_OAI21X3 U12587 ( .A(n480), .B(n481), .C(n453), .Z(n5556) );
  HS65_LL_OAI21X3 U12588 ( .A(n263), .B(n264), .C(n236), .Z(n5534) );
  HS65_LL_OAI21X3 U12589 ( .A(n305), .B(n306), .C(n278), .Z(n7148) );
  HS65_LL_OAI21X3 U12590 ( .A(n689), .B(n697), .C(n674), .Z(n5811) );
  HS65_LL_OAI21X3 U12591 ( .A(n513), .B(n521), .C(n498), .Z(n7403) );
  HS65_LL_OAI21X3 U12592 ( .A(n86), .B(n78), .C(n59), .Z(n7126) );
  HS65_LL_OAI21X3 U12593 ( .A(n170), .B(n163), .C(n155), .Z(n3284) );
  HS65_LL_OAI21X3 U12594 ( .A(n605), .B(n615), .C(n591), .Z(n8419) );
  HS65_LL_OAI21X3 U12595 ( .A(n125), .B(n135), .C(n111), .Z(n8471) );
  HS65_LL_IVX9 U12596 ( .A(n2651), .Z(n187) );
  HS65_LL_OAI21X3 U12597 ( .A(n398), .B(n392), .C(n373), .Z(n8651) );
  HS65_LL_OAI21X3 U12598 ( .A(n303), .B(n300), .C(n279), .Z(n6585) );
  HS65_LL_OAI21X3 U12599 ( .A(n85), .B(n73), .C(n58), .Z(n6473) );
  HS65_LL_OAI21X3 U12600 ( .A(n261), .B(n258), .C(n237), .Z(n4880) );
  HS65_LL_OAI21X3 U12601 ( .A(n478), .B(n475), .C(n454), .Z(n4992) );
  HS65_LL_OAI21X3 U12602 ( .A(n516), .B(n508), .C(n497), .Z(n6459) );
  HS65_LL_OAI21X3 U12603 ( .A(n692), .B(n684), .C(n673), .Z(n4866) );
  HS65_LL_OAI21X3 U12604 ( .A(n350), .B(n353), .C(n324), .Z(n8368) );
  HS65_LL_OAI21X3 U12605 ( .A(n770), .B(n758), .C(n789), .Z(n1955) );
  HS65_LL_OAI21X3 U12606 ( .A(n758), .B(n773), .C(n786), .Z(n1899) );
  HS65_LL_OAI21X3 U12607 ( .A(n881), .B(n896), .C(n909), .Z(n2275) );
  HS65_LL_OAI21X3 U12608 ( .A(n212), .B(n214), .C(n189), .Z(n4063) );
  HS65_LL_NAND2X7 U12609 ( .A(n350), .B(n328), .Z(n8607) );
  HS65_LL_OAI21X3 U12610 ( .A(n893), .B(n881), .C(n912), .Z(n2331) );
  HS65_LL_OAI21X3 U12611 ( .A(n852), .B(n840), .C(n871), .Z(n1203) );
  HS65_LL_OAI21X3 U12612 ( .A(n811), .B(n799), .C(n830), .Z(n1579) );
  HS65_LL_OAI21X3 U12613 ( .A(n124), .B(n132), .C(n112), .Z(n9079) );
  HS65_LL_OAI21X3 U12614 ( .A(n604), .B(n612), .C(n592), .Z(n9021) );
  HS65_LL_OAI21X3 U12615 ( .A(n443), .B(n429), .C(n420), .Z(n2996) );
  HS65_LL_OAI21X3 U12616 ( .A(n218), .B(n210), .C(n188), .Z(n2858) );
  HS65_LL_OAI21X3 U12617 ( .A(n437), .B(n443), .C(n407), .Z(n3410) );
  HS65_LL_OAI21X3 U12618 ( .A(n428), .B(n438), .C(n422), .Z(n4301) );
  HS65_LL_OAI21X3 U12619 ( .A(n658), .B(n655), .C(n634), .Z(n4000) );
  HS65_LL_OAI21X3 U12620 ( .A(n654), .B(n652), .C(n626), .Z(n3297) );
  HS65_LL_OAI21X3 U12621 ( .A(n34), .B(n42), .C(n19), .Z(n5749) );
  HS65_LL_OAI21X3 U12622 ( .A(n556), .B(n564), .C(n541), .Z(n7341) );
  HS65_LL_OAI21X3 U12623 ( .A(n353), .B(n341), .C(n322), .Z(n7950) );
  HS65_LL_OAI21X3 U12624 ( .A(n209), .B(n214), .C(n195), .Z(n3930) );
  HS65_LL_OAI21X3 U12625 ( .A(n215), .B(n218), .C(n200), .Z(n3065) );
  HS65_LL_OAI21X3 U12626 ( .A(n149), .B(n147), .C(n177), .Z(n4123) );
  HS65_LL_AOI12X2 U12627 ( .A(n366), .B(n8110), .C(n8111), .Z(n8109) );
  HS65_LL_OAI21X3 U12628 ( .A(n395), .B(n391), .C(n366), .Z(n7849) );
  HS65_LL_OAI21X3 U12629 ( .A(n427), .B(n438), .C(n416), .Z(n4043) );
  HS65_LL_NAND2X7 U12630 ( .A(n170), .B(n151), .Z(n3614) );
  HS65_LL_OAI21X3 U12631 ( .A(n652), .B(n660), .C(n638), .Z(n2971) );
  HS65_LL_OAI21X3 U12632 ( .A(n163), .B(n173), .C(n142), .Z(n2916) );
  HS65_LL_OAI21X3 U12633 ( .A(n655), .B(n649), .C(n636), .Z(n4263) );
  HS65_LL_OAI21X3 U12634 ( .A(n34), .B(n5478), .C(n18), .Z(n5755) );
  HS65_LL_OAI21X3 U12635 ( .A(n556), .B(n7070), .C(n540), .Z(n7347) );
  HS65_LL_OAI21X3 U12636 ( .A(n399), .B(n395), .C(n371), .Z(n8121) );
  HS65_LL_OAI21X3 U12637 ( .A(n262), .B(n256), .C(n244), .Z(n5829) );
  HS65_LL_OAI21X3 U12638 ( .A(n479), .B(n473), .C(n461), .Z(n5888) );
  HS65_LL_OAI21X3 U12639 ( .A(n691), .B(n686), .C(n670), .Z(n5680) );
  HS65_LL_OAI21X3 U12640 ( .A(n84), .B(n74), .C(n55), .Z(n7421) );
  HS65_LL_OAI21X3 U12641 ( .A(n304), .B(n298), .C(n286), .Z(n7480) );
  HS65_LL_OAI21X3 U12642 ( .A(n515), .B(n510), .C(n494), .Z(n7272) );
  HS65_LL_OAI21X3 U12643 ( .A(n214), .B(n220), .C(n193), .Z(n4070) );
  HS65_LL_OAI21X3 U12644 ( .A(n438), .B(n440), .C(n418), .Z(n4322) );
  HS65_LL_NAND2X7 U12645 ( .A(n146), .B(n177), .Z(n3624) );
  HS65_LL_OAI21X3 U12646 ( .A(n612), .B(n7700), .C(n592), .Z(n8149) );
  HS65_LL_OAI21X3 U12647 ( .A(n132), .B(n7738), .C(n112), .Z(n8172) );
  HS65_LL_NAND2X7 U12648 ( .A(n35), .B(n25), .Z(n4720) );
  HS65_LL_NAND2X7 U12649 ( .A(n557), .B(n547), .Z(n6313) );
  HS65_LL_IVX9 U12650 ( .A(n2896), .Z(n140) );
  HS65_LL_OAI21X3 U12651 ( .A(n124), .B(n7880), .C(n111), .Z(n7878) );
  HS65_LL_OAI21X3 U12652 ( .A(n604), .B(n7841), .C(n591), .Z(n7839) );
  HS65_LL_AOI12X2 U12653 ( .A(n437), .B(n416), .C(n3795), .Z(n3794) );
  HS65_LL_AOI12X2 U12654 ( .A(n215), .B(n195), .C(n3437), .Z(n3436) );
  HS65_LL_AOI12X2 U12655 ( .A(n638), .B(n3330), .C(n3331), .Z(n3329) );
  HS65_LL_NAND2X7 U12656 ( .A(n166), .B(n151), .Z(n3618) );
  HS65_LL_NAND4ABX3 U12657 ( .A(n3906), .B(n3907), .C(n3908), .D(n3909), .Z(
        n3905) );
  HS65_LL_AOI212X4 U12658 ( .A(n147), .B(n178), .C(n179), .D(n143), .E(n3910), 
        .Z(n3909) );
  HS65_LL_NAND2X7 U12659 ( .A(n461), .B(n477), .Z(n5395) );
  HS65_LL_NAND2X7 U12660 ( .A(n670), .B(n690), .Z(n5163) );
  HS65_LL_NAND2X7 U12661 ( .A(n494), .B(n514), .Z(n6755) );
  HS65_LL_AOI12X2 U12662 ( .A(n153), .B(n177), .C(n3635), .Z(n3634) );
  HS65_LL_NAND2X7 U12663 ( .A(n145), .B(n177), .Z(n3628) );
  HS65_LL_NAND2X7 U12664 ( .A(n221), .B(n202), .Z(n3521) );
  HS65_LL_AOI12X2 U12665 ( .A(n503), .B(n523), .C(n6762), .Z(n6761) );
  HS65_LL_AOI12X2 U12666 ( .A(n679), .B(n699), .C(n5170), .Z(n5169) );
  HS65_LL_AOI12X2 U12667 ( .A(n234), .B(n255), .C(n4463), .Z(n5286) );
  HS65_LL_AOI12X2 U12668 ( .A(n451), .B(n472), .C(n4502), .Z(n5401) );
  HS65_LL_AOI12X2 U12669 ( .A(n276), .B(n297), .C(n6095), .Z(n6993) );
  HS65_LL_NAND2X7 U12670 ( .A(n170), .B(n145), .Z(n3247) );
  HS65_LL_NAND3AX6 U12671 ( .A(n3187), .B(n3188), .C(n3189), .Z(n3172) );
  HS65_LL_OAI21X3 U12672 ( .A(n430), .B(n3190), .C(n405), .Z(n3189) );
  HS65_LL_NOR3AX2 U12673 ( .A(n4583), .B(n4741), .C(n4742), .Z(n4722) );
  HS65_LL_IVX9 U12674 ( .A(n3776), .Z(n410) );
  HS65_LL_NOR3AX2 U12675 ( .A(n3777), .B(n3778), .C(n3779), .Z(n3776) );
  HS65_LL_OAI21X3 U12676 ( .A(n458), .B(n462), .C(n476), .Z(n4505) );
  HS65_LL_OAI21X3 U12677 ( .A(n241), .B(n245), .C(n259), .Z(n4466) );
  HS65_LL_OAI21X3 U12678 ( .A(n283), .B(n287), .C(n301), .Z(n6098) );
  HS65_LL_OAI21X3 U12679 ( .A(n669), .B(n665), .C(n685), .Z(n5818) );
  HS65_LL_OAI21X3 U12680 ( .A(n493), .B(n489), .C(n509), .Z(n7410) );
  HS65_LL_OAI21X3 U12681 ( .A(n57), .B(n69), .C(n77), .Z(n6059) );
  HS65_LL_NAND2X7 U12682 ( .A(n212), .B(n202), .Z(n3520) );
  HS65_LL_OAI21X3 U12683 ( .A(n172), .B(n168), .C(n150), .Z(n3983) );
  HS65_LL_OAI21X3 U12684 ( .A(n561), .B(n558), .C(n538), .Z(n7095) );
  HS65_LL_OAI21X3 U12685 ( .A(n39), .B(n36), .C(n16), .Z(n5503) );
  HS65_LL_NOR3AX2 U12686 ( .A(n7937), .B(n8042), .C(n8043), .Z(n8023) );
  HS65_LL_AOI12X2 U12687 ( .A(n142), .B(n3257), .C(n3258), .Z(n3256) );
  HS65_LL_NAND2X7 U12688 ( .A(n341), .B(n317), .Z(n8340) );
  HS65_LL_NOR3AX2 U12689 ( .A(n7855), .B(n7974), .C(n7975), .Z(n7955) );
  HS65_LL_OAI21X3 U12690 ( .A(n759), .B(n1875), .C(n789), .Z(n1873) );
  HS65_LL_NOR3AX2 U12691 ( .A(n2863), .B(n3071), .C(n2944), .Z(n3055) );
  HS65_LL_OAI21X3 U12692 ( .A(n841), .B(n1123), .C(n871), .Z(n1121) );
  HS65_LL_OAI21X3 U12693 ( .A(n800), .B(n1499), .C(n830), .Z(n1497) );
  HS65_LL_OAI21X3 U12694 ( .A(n882), .B(n2251), .C(n912), .Z(n2249) );
  HS65_LL_OAI21X3 U12695 ( .A(n169), .B(n180), .C(n145), .Z(n3052) );
  HS65_LL_NAND2X7 U12696 ( .A(n610), .B(n593), .Z(n7625) );
  HS65_LL_NAND2X7 U12697 ( .A(n130), .B(n113), .Z(n7665) );
  HS65_LL_NOR4ABX2 U12698 ( .A(n5473), .B(n5474), .C(n5475), .D(n5476), .Z(
        n5467) );
  HS65_LL_AOI212X4 U12699 ( .A(n45), .B(n14), .C(n10), .D(n46), .E(n5477), .Z(
        n5474) );
  HS65_LL_NOR4ABX2 U12700 ( .A(n7065), .B(n7066), .C(n7067), .D(n7068), .Z(
        n7059) );
  HS65_LL_AOI212X4 U12701 ( .A(n567), .B(n536), .C(n532), .D(n568), .E(n7069), 
        .Z(n7066) );
  HS65_LL_AOI12X2 U12702 ( .A(n330), .B(n347), .C(n8574), .Z(n8573) );
  HS65_LL_OAI21X3 U12703 ( .A(n607), .B(n602), .C(n582), .Z(n8136) );
  HS65_LL_OAI21X3 U12704 ( .A(n127), .B(n122), .C(n102), .Z(n8187) );
  HS65_LL_OAI21X3 U12705 ( .A(n147), .B(n142), .C(n164), .Z(n4163) );
  HS65_LL_OAI21X3 U12706 ( .A(n167), .B(n3912), .C(n155), .Z(n4162) );
  HS65_LL_OAI21X3 U12707 ( .A(n563), .B(n558), .C(n532), .Z(n7255) );
  HS65_LL_OAI21X3 U12708 ( .A(n41), .B(n36), .C(n10), .Z(n5663) );
  HS65_LL_NAND2X7 U12709 ( .A(n334), .B(n352), .Z(n8602) );
  HS65_LL_OAI21X3 U12710 ( .A(n439), .B(n2843), .C(n407), .Z(n2841) );
  HS65_LL_AOI12X2 U12711 ( .A(n462), .B(n4980), .C(n4981), .Z(n4979) );
  HS65_LL_AOI12X2 U12712 ( .A(n287), .B(n6573), .C(n6574), .Z(n6572) );
  HS65_LL_AOI12X2 U12713 ( .A(n489), .B(n6447), .C(n6448), .Z(n6446) );
  HS65_LL_AOI12X2 U12714 ( .A(n665), .B(n4854), .C(n4855), .Z(n4853) );
  HS65_LL_OAI21X3 U12715 ( .A(n656), .B(n2895), .C(n626), .Z(n2893) );
  HS65_LL_OAI21X3 U12716 ( .A(n213), .B(n3897), .C(n200), .Z(n4224) );
  HS65_LL_NAND2X7 U12717 ( .A(n407), .B(n433), .Z(n3831) );
  HS65_LL_AOI12X2 U12718 ( .A(n584), .B(n7830), .C(n8400), .Z(n8399) );
  HS65_LL_AOI12X2 U12719 ( .A(n104), .B(n7928), .C(n8452), .Z(n8451) );
  HS65_LL_NAND2X7 U12720 ( .A(n200), .B(n224), .Z(n3476) );
  HS65_LL_NOR4ABX2 U12721 ( .A(n3908), .B(n3985), .C(n3986), .D(n3987), .Z(
        n3979) );
  HS65_LL_AOI212X4 U12722 ( .A(n169), .B(n143), .C(n142), .D(n175), .E(n3988), 
        .Z(n3985) );
  HS65_LL_NAND2X7 U12723 ( .A(n191), .B(n220), .Z(n3495) );
  HS65_LL_NOR3AX2 U12724 ( .A(n3144), .B(n3145), .C(n2978), .Z(n3123) );
  HS65_LL_NOR3AX2 U12725 ( .A(n2943), .B(n2944), .C(n2866), .Z(n2921) );
  HS65_LL_NAND2X7 U12726 ( .A(n611), .B(n590), .Z(n7687) );
  HS65_LL_NAND2X7 U12727 ( .A(n131), .B(n110), .Z(n7725) );
  HS65_LL_OAI21X3 U12728 ( .A(n480), .B(n4506), .C(n454), .Z(n4504) );
  HS65_LL_OAI21X3 U12729 ( .A(n263), .B(n4467), .C(n237), .Z(n4465) );
  HS65_LL_OAI21X3 U12730 ( .A(n305), .B(n6099), .C(n279), .Z(n6097) );
  HS65_LL_OAI21X3 U12731 ( .A(n689), .B(n5492), .C(n673), .Z(n5817) );
  HS65_LL_OAI21X3 U12732 ( .A(n513), .B(n7084), .C(n497), .Z(n7409) );
  HS65_LL_OAI21X3 U12733 ( .A(n86), .B(n6060), .C(n58), .Z(n6058) );
  HS65_LL_NAND4ABX3 U12734 ( .A(n8255), .B(n8091), .C(n8490), .D(n8199), .Z(
        n8487) );
  HS65_LL_OAI21X3 U12735 ( .A(n397), .B(n394), .C(n369), .Z(n8490) );
  HS65_LL_NAND2X7 U12736 ( .A(n191), .B(n224), .Z(n3091) );
  HS65_LL_OAI21X3 U12737 ( .A(n417), .B(n415), .C(n435), .Z(n4306) );
  HS65_LL_NAND2X7 U12738 ( .A(n419), .B(n433), .Z(n3376) );
  HS65_LL_NAND2X7 U12739 ( .A(n96), .B(n137), .Z(n8789) );
  HS65_LL_NAND2X7 U12740 ( .A(n20), .B(n37), .Z(n5031) );
  HS65_LL_NAND2X7 U12741 ( .A(n542), .B(n559), .Z(n6624) );
  HS65_LL_OAI21X3 U12742 ( .A(n174), .B(n168), .C(n143), .Z(n4094) );
  HS65_LL_OAI21X3 U12743 ( .A(n194), .B(n192), .C(n223), .Z(n4173) );
  HS65_LL_NAND2X7 U12744 ( .A(n146), .B(n180), .Z(n3625) );
  HS65_LL_OAI21X3 U12745 ( .A(n583), .B(n584), .C(n610), .Z(n8135) );
  HS65_LL_OAI21X3 U12746 ( .A(n103), .B(n104), .C(n130), .Z(n8186) );
  HS65_LL_OAI21X3 U12747 ( .A(n640), .B(n638), .C(n659), .Z(n3138) );
  HS65_LL_NOR4ABX2 U12748 ( .A(n3607), .B(n3285), .C(n3654), .D(n3636), .Z(
        n3990) );
  HS65_LL_OAI21X3 U12749 ( .A(n333), .B(n322), .C(n356), .Z(n8618) );
  HS65_LL_OAI21X3 U12750 ( .A(n320), .B(n322), .C(n340), .Z(n8038) );
  HS65_LL_NAND2X7 U12751 ( .A(n146), .B(n167), .Z(n3026) );
  HS65_LL_NOR4ABX2 U12752 ( .A(n6820), .B(n6821), .C(n6822), .D(n6823), .Z(
        n6813) );
  HS65_LL_NOR4ABX2 U12753 ( .A(n5228), .B(n5229), .C(n5230), .D(n5231), .Z(
        n5221) );
  HS65_LL_OAI21X3 U12754 ( .A(n367), .B(n366), .C(n396), .Z(n8660) );
  HS65_LL_OAI21X3 U12755 ( .A(n260), .B(n252), .C(n246), .Z(n4738) );
  HS65_LL_OAI21X3 U12756 ( .A(n477), .B(n469), .C(n463), .Z(n4799) );
  HS65_LL_OAI21X3 U12757 ( .A(n302), .B(n294), .C(n288), .Z(n6392) );
  HS65_LL_OAI21X3 U12758 ( .A(n83), .B(n89), .C(n67), .Z(n6353) );
  HS65_LL_OAI21X3 U12759 ( .A(n514), .B(n526), .C(n492), .Z(n6246) );
  HS65_LL_OAI21X3 U12760 ( .A(n690), .B(n702), .C(n668), .Z(n4653) );
  HS65_LL_OAI21X3 U12761 ( .A(n99), .B(n104), .C(n136), .Z(n7879) );
  HS65_LL_OAI21X3 U12762 ( .A(n579), .B(n584), .C(n616), .Z(n7840) );
  HS65_LL_NOR4ABX2 U12763 ( .A(n4978), .B(n4993), .C(n5383), .D(n5403), .Z(
        n5632) );
  HS65_LL_NOR4ABX2 U12764 ( .A(n4852), .B(n4867), .C(n5151), .D(n5172), .Z(
        n5575) );
  HS65_LL_NOR4ABX2 U12765 ( .A(n6445), .B(n6460), .C(n6743), .D(n6764), .Z(
        n7167) );
  HS65_LL_NOR4ABX2 U12766 ( .A(n6571), .B(n6586), .C(n6975), .D(n6995), .Z(
        n7224) );
  HS65_LL_NOR4ABX2 U12767 ( .A(n4925), .B(n4881), .C(n5268), .D(n5288), .Z(
        n5606) );
  HS65_LL_OAI21X3 U12768 ( .A(n35), .B(n47), .C(n11), .Z(n4576) );
  HS65_LL_OAI21X3 U12769 ( .A(n557), .B(n569), .C(n533), .Z(n6169) );
  HS65_LL_NAND2X7 U12770 ( .A(n15), .B(n35), .Z(n5041) );
  HS65_LL_NAND2X7 U12771 ( .A(n537), .B(n557), .Z(n6634) );
  HS65_LL_OAI21X3 U12772 ( .A(n363), .B(n366), .C(n389), .Z(n7969) );
  HS65_LL_IVX9 U12773 ( .A(n2897), .Z(n141) );
  HS65_LL_NAND2X7 U12774 ( .A(n399), .B(n365), .Z(n8103) );
  HS65_LL_NAND2X7 U12775 ( .A(n344), .B(n322), .Z(n8572) );
  HS65_LL_NAND2X7 U12776 ( .A(n326), .B(n344), .Z(n8555) );
  HS65_LL_NAND2X7 U12777 ( .A(n215), .B(n190), .Z(n3092) );
  HS65_LL_NOR4ABX2 U12778 ( .A(n8340), .B(n8577), .C(n8366), .D(n8557), .Z(
        n8921) );
  HS65_LL_NOR3AX2 U12779 ( .A(n6151), .B(n6152), .C(n6153), .Z(n6139) );
  HS65_LL_OAI21X3 U12780 ( .A(n564), .B(n6154), .C(n541), .Z(n6151) );
  HS65_LL_NOR3AX2 U12781 ( .A(n4558), .B(n4559), .C(n4560), .Z(n4546) );
  HS65_LL_OAI21X3 U12782 ( .A(n42), .B(n4561), .C(n19), .Z(n4558) );
  HS65_LL_NOR3AX2 U12783 ( .A(n4754), .B(n4755), .C(n4756), .Z(n4744) );
  HS65_LL_OAI21X3 U12784 ( .A(n264), .B(n4757), .C(n236), .Z(n4754) );
  HS65_LL_NOR3AX2 U12785 ( .A(n6228), .B(n6229), .C(n6230), .Z(n6216) );
  HS65_LL_OAI21X3 U12786 ( .A(n521), .B(n6231), .C(n498), .Z(n6228) );
  HS65_LL_NOR3AX2 U12787 ( .A(n4781), .B(n4782), .C(n4783), .Z(n4770) );
  HS65_LL_OAI21X3 U12788 ( .A(n481), .B(n4784), .C(n453), .Z(n4781) );
  HS65_LL_NOR3AX2 U12789 ( .A(n6374), .B(n6375), .C(n6376), .Z(n6363) );
  HS65_LL_OAI21X3 U12790 ( .A(n306), .B(n6377), .C(n278), .Z(n6374) );
  HS65_LL_NOR3AX2 U12791 ( .A(n6335), .B(n6336), .C(n6337), .Z(n6324) );
  HS65_LL_OAI21X3 U12792 ( .A(n78), .B(n6338), .C(n59), .Z(n6335) );
  HS65_LL_NOR3AX2 U12793 ( .A(n4635), .B(n4636), .C(n4637), .Z(n4623) );
  HS65_LL_OAI21X3 U12794 ( .A(n697), .B(n4638), .C(n674), .Z(n4635) );
  HS65_LL_OAI21X3 U12795 ( .A(n342), .B(n352), .C(n335), .Z(n8877) );
  HS65_LL_NAND2X7 U12796 ( .A(n9), .B(n36), .Z(n5081) );
  HS65_LL_NAND2X7 U12797 ( .A(n531), .B(n558), .Z(n6674) );
  HS65_LL_NOR4ABX2 U12798 ( .A(n3099), .B(n3520), .C(n3493), .D(n3513), .Z(
        n4067) );
  HS65_LL_NOR3AX2 U12799 ( .A(n8359), .B(n8360), .C(n8361), .Z(n8350) );
  HS65_LL_OAI21X3 U12800 ( .A(n609), .B(n606), .C(n576), .Z(n7621) );
  HS65_LL_OAI21X3 U12801 ( .A(n129), .B(n126), .C(n96), .Z(n7661) );
  HS65_LL_OAI21X3 U12802 ( .A(n656), .B(n661), .C(n624), .Z(n3945) );
  HS65_LL_NAND2X7 U12803 ( .A(n406), .B(n439), .Z(n3372) );
  HS65_LL_NAND2X7 U12804 ( .A(n676), .B(n688), .Z(n5183) );
  HS65_LL_NAND2X7 U12805 ( .A(n500), .B(n512), .Z(n6775) );
  HS65_LL_NAND2X7 U12806 ( .A(n148), .B(n177), .Z(n3610) );
  HS65_LL_NOR4ABX2 U12807 ( .A(n8253), .B(n8122), .C(n8111), .D(n8270), .Z(
        n8973) );
  HS65_LL_OAI21X3 U12808 ( .A(n415), .B(n420), .C(n442), .Z(n2842) );
  HS65_LL_NAND2X7 U12809 ( .A(n625), .B(n656), .Z(n3318) );
  HS65_LL_NAND2X7 U12810 ( .A(n88), .B(n64), .Z(n6836) );
  HS65_LL_NAND2X7 U12811 ( .A(n253), .B(n233), .Z(n5244) );
  HS65_LL_NAND2X7 U12812 ( .A(n470), .B(n450), .Z(n5359) );
  HS65_LL_NAND2X7 U12813 ( .A(n700), .B(n678), .Z(n5126) );
  HS65_LL_NAND2X7 U12814 ( .A(n295), .B(n275), .Z(n6951) );
  HS65_LL_NAND2X7 U12815 ( .A(n524), .B(n502), .Z(n6718) );
  HS65_LL_OAI21X3 U12816 ( .A(n168), .B(n165), .C(n148), .Z(n4101) );
  HS65_LL_OAI21X3 U12817 ( .A(n439), .B(n430), .C(n405), .Z(n3965) );
  HS65_LL_NOR4ABX2 U12818 ( .A(n8607), .B(n8608), .C(n8609), .D(n8610), .Z(
        n8595) );
  HS65_LL_NAND2X7 U12819 ( .A(n203), .B(n213), .Z(n3087) );
  HS65_LL_NOR3AX2 U12820 ( .A(n3401), .B(n3402), .C(n3403), .Z(n3390) );
  HS65_LL_OAI21X3 U12821 ( .A(n417), .B(n3365), .C(n431), .Z(n3401) );
  HS65_LL_NOR3AX2 U12822 ( .A(n3120), .B(n3121), .C(n3122), .Z(n3107) );
  HS65_LL_OAI21X3 U12823 ( .A(n194), .B(n3080), .C(n225), .Z(n3120) );
  HS65_LL_OAI21X3 U12824 ( .A(n633), .B(n638), .C(n651), .Z(n2894) );
  HS65_LL_NAND2X7 U12825 ( .A(n375), .B(n384), .Z(n8198) );
  HS65_LL_NOR4ABX2 U12826 ( .A(n4714), .B(n5051), .C(n4664), .D(n5030), .Z(
        n5511) );
  HS65_LL_NOR4ABX2 U12827 ( .A(n6307), .B(n6644), .C(n6257), .D(n6623), .Z(
        n7103) );
  HS65_LL_OAI21X3 U12828 ( .A(n126), .B(n137), .C(n98), .Z(n9097) );
  HS65_LL_OAI21X3 U12829 ( .A(n606), .B(n617), .C(n578), .Z(n9039) );
  HS65_LL_NAND2X7 U12830 ( .A(n665), .B(n692), .Z(n5204) );
  HS65_LL_NAND2X7 U12831 ( .A(n489), .B(n516), .Z(n6796) );
  HS65_LL_NAND2X7 U12832 ( .A(n107), .B(n125), .Z(n7912) );
  HS65_LL_NAND2X7 U12833 ( .A(n587), .B(n605), .Z(n7814) );
  HS65_LL_IVX9 U12834 ( .A(n2755), .Z(n361) );
  HS65_LL_OAI21X3 U12835 ( .A(n422), .B(n420), .C(n428), .Z(n3201) );
  HS65_LL_NOR4ABX2 U12836 ( .A(n7790), .B(n7693), .C(n8151), .D(n8152), .Z(
        n8142) );
  HS65_LL_NOR4ABX2 U12837 ( .A(n7889), .B(n7731), .C(n8174), .D(n8175), .Z(
        n8165) );
  HS65_LL_NAND2X7 U12838 ( .A(n370), .B(n397), .Z(n8221) );
  HS65_LL_NAND2X7 U12839 ( .A(n147), .B(n167), .Z(n3272) );
  HS65_LL_NAND2X7 U12840 ( .A(n654), .B(n630), .Z(n3673) );
  HS65_LL_OAI21X3 U12841 ( .A(n326), .B(n322), .C(n351), .Z(n8358) );
  HS65_LL_NOR3AX2 U12842 ( .A(n3275), .B(n3276), .C(n3277), .Z(n3263) );
  HS65_LL_OAI21X3 U12843 ( .A(n149), .B(n3236), .C(n179), .Z(n3275) );
  HS65_LL_NOR4ABX2 U12844 ( .A(n3382), .B(n3874), .C(n3848), .D(n3867), .Z(
        n4319) );
  HS65_LL_OAI21X3 U12845 ( .A(n234), .B(n4897), .C(n258), .Z(n4905) );
  HS65_LL_OAI21X3 U12846 ( .A(n451), .B(n4950), .C(n475), .Z(n4958) );
  HS65_LL_OAI21X3 U12847 ( .A(n276), .B(n6543), .C(n300), .Z(n6551) );
  HS65_LL_OAI21X3 U12848 ( .A(n63), .B(n6490), .C(n73), .Z(n6498) );
  HS65_LL_OAI21X3 U12849 ( .A(n503), .B(n6415), .C(n508), .Z(n6423) );
  HS65_LL_OAI21X3 U12850 ( .A(n679), .B(n4822), .C(n684), .Z(n4830) );
  HS65_LL_NAND2X7 U12851 ( .A(n556), .B(n543), .Z(n6644) );
  HS65_LL_NAND2X7 U12852 ( .A(n34), .B(n21), .Z(n5051) );
  HS65_LL_OAI21X3 U12853 ( .A(n203), .B(n188), .C(n216), .Z(n3113) );
  HS65_LL_OAI21X3 U12854 ( .A(n609), .B(n614), .C(n580), .Z(n8416) );
  HS65_LL_OAI21X3 U12855 ( .A(n129), .B(n134), .C(n100), .Z(n8468) );
  HS65_LL_NAND2X7 U12856 ( .A(n438), .B(n409), .Z(n3800) );
  HS65_LL_NOR3AX2 U12857 ( .A(n7987), .B(n7988), .C(n7989), .Z(n7977) );
  HS65_LL_OAI21X3 U12858 ( .A(n392), .B(n7743), .C(n373), .Z(n7987) );
  HS65_LL_NAND2X7 U12859 ( .A(n437), .B(n412), .Z(n3788) );
  HS65_LL_NAND2X7 U12860 ( .A(n103), .B(n131), .Z(n8446) );
  HS65_LL_NAND2X7 U12861 ( .A(n583), .B(n611), .Z(n8394) );
  HS65_LL_NAND2X7 U12862 ( .A(n172), .B(n143), .Z(n3606) );
  HS65_LL_NAND2X7 U12863 ( .A(n173), .B(n143), .Z(n3248) );
  HS65_LL_OAI21X3 U12864 ( .A(n172), .B(n166), .C(n149), .Z(n3281) );
  HS65_LL_OAI21X3 U12865 ( .A(n888), .B(n885), .C(n914), .Z(n2328) );
  HS65_LL_OAI21X3 U12866 ( .A(n342), .B(n355), .C(n334), .Z(n8364) );
  HS65_LL_OAI21X3 U12867 ( .A(n765), .B(n762), .C(n791), .Z(n1952) );
  HS65_LL_NAND2X7 U12868 ( .A(n19), .B(n40), .Z(n5038) );
  HS65_LL_NAND2X7 U12869 ( .A(n541), .B(n562), .Z(n6631) );
  HS65_LL_NAND2X7 U12870 ( .A(n453), .B(n482), .Z(n5392) );
  HS65_LL_NAND2X7 U12871 ( .A(n674), .B(n695), .Z(n5160) );
  HS65_LL_NAND2X7 U12872 ( .A(n278), .B(n307), .Z(n6984) );
  HS65_LL_NAND2X7 U12873 ( .A(n498), .B(n519), .Z(n6752) );
  HS65_LL_OAI21X3 U12874 ( .A(n847), .B(n844), .C(n873), .Z(n1200) );
  HS65_LL_OAI21X3 U12875 ( .A(n806), .B(n803), .C(n832), .Z(n1576) );
  HS65_LL_NAND2X7 U12876 ( .A(n478), .B(n452), .Z(n5462) );
  HS65_LL_NAND2X7 U12877 ( .A(n692), .B(n680), .Z(n5232) );
  HS65_LL_NAND2X7 U12878 ( .A(n516), .B(n504), .Z(n6824) );
  HS65_LL_OAI21X3 U12879 ( .A(n39), .B(n33), .C(n17), .Z(n4662) );
  HS65_LL_OAI21X3 U12880 ( .A(n561), .B(n555), .C(n539), .Z(n6255) );
  HS65_LL_NAND3AX6 U12881 ( .A(n7691), .B(n7692), .C(n7693), .Z(n7689) );
  HS65_LL_NAND3AX6 U12882 ( .A(n7729), .B(n7730), .C(n7731), .Z(n7727) );
  HS65_LL_OAI21X3 U12883 ( .A(n209), .B(n221), .C(n194), .Z(n3062) );
  HS65_LL_OAI21X3 U12884 ( .A(n390), .B(n393), .C(n370), .Z(n8118) );
  HS65_LL_OAI21X3 U12885 ( .A(n326), .B(n325), .C(n342), .Z(n8050) );
  HS65_LL_OAI21X3 U12886 ( .A(n372), .B(n374), .C(n390), .Z(n7982) );
  HS65_LL_OAI21X3 U12887 ( .A(n658), .B(n650), .C(n635), .Z(n3294) );
  HS65_LL_OAI21X3 U12888 ( .A(n310), .B(n299), .C(n285), .Z(n6582) );
  HS65_LL_OAI21X3 U12889 ( .A(n82), .B(n76), .C(n56), .Z(n6470) );
  HS65_LL_OAI21X3 U12890 ( .A(n268), .B(n257), .C(n243), .Z(n4877) );
  HS65_LL_OAI21X3 U12891 ( .A(n485), .B(n474), .C(n460), .Z(n4989) );
  HS65_LL_OAI21X3 U12892 ( .A(n518), .B(n512), .C(n496), .Z(n6456) );
  HS65_LL_OAI21X3 U12893 ( .A(n694), .B(n688), .C(n672), .Z(n4863) );
  HS65_LL_NAND2X7 U12894 ( .A(n10), .B(n40), .Z(n4706) );
  HS65_LL_NAND2X7 U12895 ( .A(n532), .B(n562), .Z(n6299) );
  HS65_LL_NAND2X7 U12896 ( .A(n464), .B(n482), .Z(n4972) );
  HS65_LL_NAND2X7 U12897 ( .A(n666), .B(n695), .Z(n4844) );
  HS65_LL_NAND2X7 U12898 ( .A(n490), .B(n519), .Z(n6437) );
  HS65_LL_OAI21X3 U12899 ( .A(n427), .B(n441), .C(n417), .Z(n3407) );
  HS65_LL_OAI21X3 U12900 ( .A(n631), .B(n3311), .C(n652), .Z(n3308) );
  HS65_LL_OAI21X3 U12901 ( .A(n378), .B(n8080), .C(n395), .Z(n8089) );
  HS65_LL_OAI21X3 U12902 ( .A(n330), .B(n8324), .C(n353), .Z(n8321) );
  HS65_LL_NAND2X7 U12903 ( .A(n221), .B(n196), .Z(n3490) );
  HS65_LL_NAND2X7 U12904 ( .A(n191), .B(n213), .Z(n2953) );
  HS65_LL_NAND2X7 U12905 ( .A(n419), .B(n439), .Z(n3180) );
  HS65_LL_NAND2X7 U12906 ( .A(n637), .B(n656), .Z(n3154) );
  HS65_LL_OAI21X3 U12907 ( .A(n585), .B(n8385), .C(n615), .Z(n8382) );
  HS65_LL_OAI21X3 U12908 ( .A(n105), .B(n8437), .C(n135), .Z(n8434) );
  HS65_LL_NAND2X7 U12909 ( .A(n533), .B(n556), .Z(n6155) );
  HS65_LL_NAND2X7 U12910 ( .A(n11), .B(n34), .Z(n4562) );
  HS65_LL_NAND2X7 U12911 ( .A(n216), .B(n196), .Z(n3452) );
  HS65_LL_OAI21X3 U12912 ( .A(n24), .B(n4683), .C(n29), .Z(n4692) );
  HS65_LL_OAI21X3 U12913 ( .A(n546), .B(n6276), .C(n551), .Z(n6285) );
  HS65_LL_OAI21X3 U12914 ( .A(n413), .B(n3365), .C(n443), .Z(n3362) );
  HS65_LL_OAI21X3 U12915 ( .A(n198), .B(n3080), .C(n218), .Z(n3077) );
  HS65_LL_NAND2X7 U12916 ( .A(n436), .B(n409), .Z(n3809) );
  HS65_LL_NAND2X7 U12917 ( .A(n33), .B(n22), .Z(n5018) );
  HS65_LL_NAND2X7 U12918 ( .A(n555), .B(n544), .Z(n6611) );
  HS65_LL_NAND2X7 U12919 ( .A(n147), .B(n165), .Z(n3607) );
  HS65_LL_NAND2X7 U12920 ( .A(n637), .B(n650), .Z(n3323) );
  HS65_LL_NAND2X7 U12921 ( .A(n327), .B(n345), .Z(n8501) );
  HS65_LL_OAI21X3 U12922 ( .A(n542), .B(n543), .C(n561), .Z(n6146) );
  HS65_LL_OAI21X3 U12923 ( .A(n20), .B(n21), .C(n39), .Z(n4553) );
  HS65_LL_NAND2X7 U12924 ( .A(n419), .B(n441), .Z(n3377) );
  HS65_LL_NAND2X7 U12925 ( .A(n411), .B(n432), .Z(n3777) );
  HS65_LL_OAI21X3 U12926 ( .A(n406), .B(n408), .C(n427), .Z(n3186) );
  HS65_LL_OAI21X3 U12927 ( .A(n203), .B(n202), .C(n209), .Z(n2959) );
  HS65_LL_OAI21X3 U12928 ( .A(n238), .B(n240), .C(n268), .Z(n4749) );
  HS65_LL_OAI21X3 U12929 ( .A(n499), .B(n500), .C(n518), .Z(n6223) );
  HS65_LL_OAI21X3 U12930 ( .A(n455), .B(n457), .C(n485), .Z(n4776) );
  HS65_LL_OAI21X3 U12931 ( .A(n280), .B(n282), .C(n310), .Z(n6369) );
  HS65_LL_OAI21X3 U12932 ( .A(n60), .B(n62), .C(n82), .Z(n6330) );
  HS65_LL_OAI21X3 U12933 ( .A(n675), .B(n676), .C(n694), .Z(n4630) );
  HS65_LL_OAI21X3 U12934 ( .A(n625), .B(n627), .C(n658), .Z(n3159) );
  HS65_LL_OAI21X3 U12935 ( .A(n153), .B(n3236), .C(n163), .Z(n3233) );
  HS65_LL_NAND2X7 U12936 ( .A(n110), .B(n122), .Z(n8778) );
  HS65_LL_NAND2X7 U12937 ( .A(n590), .B(n602), .Z(n8688) );
  HS65_LL_NAND2X7 U12938 ( .A(n457), .B(n469), .Z(n5381) );
  HS65_LL_NAND2X7 U12939 ( .A(n240), .B(n252), .Z(n5266) );
  HS65_LL_NAND2X7 U12940 ( .A(n282), .B(n294), .Z(n6973) );
  HS65_LL_NAND2X7 U12941 ( .A(n676), .B(n702), .Z(n5149) );
  HS65_LL_NAND2X7 U12942 ( .A(n500), .B(n526), .Z(n6741) );
  HS65_LL_NAND2X7 U12943 ( .A(n62), .B(n89), .Z(n6858) );
  HS65_LL_OAI21X3 U12944 ( .A(n158), .B(n142), .C(n169), .Z(n3268) );
  HS65_LL_AOI12X2 U12945 ( .A(n605), .B(n576), .C(n8726), .Z(n8723) );
  HS65_LL_AOI12X2 U12946 ( .A(n125), .B(n96), .C(n8816), .Z(n8813) );
  HS65_LL_NAND2X7 U12947 ( .A(n694), .B(n666), .Z(n5140) );
  HS65_LL_NOR2X6 U12948 ( .A(n351), .B(n354), .Z(n8362) );
  HS65_LL_NAND2X7 U12949 ( .A(n146), .B(n173), .Z(n3243) );
  HS65_LL_NAND2X7 U12950 ( .A(n21), .B(n47), .Z(n5027) );
  HS65_LL_NAND2X7 U12951 ( .A(n543), .B(n569), .Z(n6620) );
  HS65_LL_OAI21X3 U12952 ( .A(n406), .B(n420), .C(n436), .Z(n3395) );
  HS65_LL_OAI21X3 U12953 ( .A(n280), .B(n287), .C(n302), .Z(n6545) );
  HS65_LL_OAI21X3 U12954 ( .A(n60), .B(n69), .C(n83), .Z(n6492) );
  HS65_LL_OAI21X3 U12955 ( .A(n238), .B(n245), .C(n260), .Z(n4899) );
  HS65_LL_OAI21X3 U12956 ( .A(n455), .B(n462), .C(n477), .Z(n4952) );
  HS65_LL_OAI21X3 U12957 ( .A(n499), .B(n489), .C(n514), .Z(n6417) );
  HS65_LL_OAI21X3 U12958 ( .A(n675), .B(n665), .C(n690), .Z(n4824) );
  HS65_LL_NAND2X7 U12959 ( .A(n107), .B(n119), .Z(n8819) );
  HS65_LL_NAND2X7 U12960 ( .A(n587), .B(n599), .Z(n8729) );
  HS65_LL_BFX9 U12961 ( .A(n9149), .Z(n9145) );
  HS65_LL_NOR2X6 U12962 ( .A(n376), .B(n374), .Z(n8301) );
  HS65_LL_NOR2X6 U12963 ( .A(n889), .B(n890), .Z(n2325) );
  HS65_LL_NOR2X6 U12964 ( .A(n766), .B(n767), .Z(n1949) );
  HS65_LL_NOR2X6 U12965 ( .A(n848), .B(n849), .Z(n1197) );
  HS65_LL_NOR2X6 U12966 ( .A(n807), .B(n808), .Z(n1573) );
  HS65_LL_NAND2X7 U12967 ( .A(n105), .B(n123), .Z(n7925) );
  HS65_LL_NAND2X7 U12968 ( .A(n585), .B(n603), .Z(n7827) );
  HS65_LL_NOR2X6 U12969 ( .A(n653), .B(n649), .Z(n3291) );
  HS65_LL_NOR2X6 U12970 ( .A(n302), .B(n298), .Z(n6579) );
  HS65_LL_NOR2X6 U12971 ( .A(n83), .B(n74), .Z(n6467) );
  HS65_LL_NOR2X6 U12972 ( .A(n260), .B(n256), .Z(n4874) );
  HS65_LL_NOR2X6 U12973 ( .A(n477), .B(n473), .Z(n4986) );
  HS65_LL_NOR2X6 U12974 ( .A(n514), .B(n510), .Z(n6453) );
  HS65_LL_NOR2X6 U12975 ( .A(n690), .B(n686), .Z(n4860) );
  HS65_LL_NOR2X6 U12976 ( .A(n216), .B(n220), .Z(n3059) );
  HS65_LL_NOR2X6 U12977 ( .A(n436), .B(n440), .Z(n3404) );
  HS65_LLS_XNOR2X6 U12978 ( .A(n2638), .B(n2644), .Z(n2690) );
  HS65_LLS_XNOR2X6 U12979 ( .A(n2692), .B(n2634), .Z(n2643) );
  HS65_LL_NOR2X6 U12980 ( .A(n35), .B(n31), .Z(n4659) );
  HS65_LL_NOR2X6 U12981 ( .A(n557), .B(n553), .Z(n6252) );
  HS65_LL_BFX9 U12982 ( .A(n9149), .Z(n9143) );
  HS65_LL_BFX9 U12983 ( .A(n9149), .Z(n9144) );
  HS65_LL_NAND3AX6 U12984 ( .A(n3662), .B(n3663), .C(n3664), .Z(n3661) );
  HS65_LL_NAND3AX6 U12985 ( .A(n3419), .B(n3420), .C(n3421), .Z(n3418) );
  HS65_LL_NAND3AX6 U12986 ( .A(n3543), .B(n3544), .C(n3545), .Z(n3542) );
  HS65_LL_BFX9 U12987 ( .A(n9134), .Z(n9129) );
  HS65_LL_BFX9 U12988 ( .A(n9134), .Z(n9130) );
  HS65_LL_OAI21X3 U12989 ( .A(n593), .B(n590), .C(n609), .Z(n8147) );
  HS65_LL_OAI21X3 U12990 ( .A(n113), .B(n110), .C(n129), .Z(n8170) );
  HS65_LL_BFX9 U12991 ( .A(n9133), .Z(n9131) );
  HS65_LL_OAI21X3 U12992 ( .A(n625), .B(n638), .C(n653), .Z(n3341) );
  HS65_LL_NAND3AX6 U12993 ( .A(n5002), .B(n5003), .C(n5004), .Z(n5001) );
  HS65_LL_NAND3AX6 U12994 ( .A(n6595), .B(n6596), .C(n6597), .Z(n6594) );
  HS65_LL_NAND2X7 U12995 ( .A(n653), .B(n628), .Z(n3694) );
  HS65_LL_NAND2X7 U12996 ( .A(n377), .B(n400), .Z(n8304) );
  HS65_LL_OAI21X3 U12997 ( .A(n580), .B(n8385), .C(n603), .Z(n8410) );
  HS65_LL_OAI21X3 U12998 ( .A(n100), .B(n8437), .C(n123), .Z(n8462) );
  HS65_LL_NAND2X7 U12999 ( .A(n408), .B(n432), .Z(n3837) );
  HS65_LL_NAND2X7 U13000 ( .A(n202), .B(n226), .Z(n3482) );
  HS65_LL_NAND2X7 U13001 ( .A(n607), .B(n579), .Z(n7688) );
  HS65_LL_NAND2X7 U13002 ( .A(n127), .B(n99), .Z(n7726) );
  HS65_LL_NOR2X6 U13003 ( .A(n629), .B(n628), .Z(n3340) );
  HS65_LL_NOR2X6 U13004 ( .A(n197), .B(n196), .Z(n3111) );
  HS65_LL_NOR2X6 U13005 ( .A(n152), .B(n151), .Z(n3267) );
  HS65_LL_NOR2X6 U13006 ( .A(n169), .B(n165), .Z(n3278) );
  HS65_LL_NAND3AX6 U13007 ( .A(n8500), .B(n8501), .C(n8502), .Z(n8499) );
  HS65_LL_NOR2X6 U13008 ( .A(n607), .B(n617), .Z(n8415) );
  HS65_LL_NOR2X6 U13009 ( .A(n127), .B(n137), .Z(n8467) );
  HS65_LL_NOR2X6 U13010 ( .A(n195), .B(n3417), .Z(n3489) );
  HS65_LL_NOR2X6 U13011 ( .A(n495), .B(n6714), .Z(n6739) );
  HS65_LL_NOR2X6 U13012 ( .A(n671), .B(n5122), .Z(n5147) );
  HS65_LL_NOR2X6 U13013 ( .A(n459), .B(n5355), .Z(n5379) );
  HS65_LL_NOR2X6 U13014 ( .A(n284), .B(n6947), .Z(n6971) );
  HS65_LL_AOI12X2 U13015 ( .A(n350), .B(n335), .C(n8606), .Z(n8603) );
  HS65_LL_NOR3AX2 U13016 ( .A(n6150), .B(n535), .C(n6614), .Z(n7248) );
  HS65_LL_IVX9 U13017 ( .A(n6630), .Z(n535) );
  HS65_LL_NOR3AX2 U13018 ( .A(n4557), .B(n13), .C(n5021), .Z(n5656) );
  HS65_LL_IVX9 U13019 ( .A(n5037), .Z(n13) );
  HS65_LL_MX41X7 U13020 ( .D0(n578), .S0(n610), .D1(n600), .S1(n592), .D2(n615), .S2(n580), .D3(n604), .S3(n591), .Z(n8724) );
  HS65_LL_MX41X7 U13021 ( .D0(n98), .S0(n130), .D1(n120), .S1(n112), .D2(n135), 
        .S2(n100), .D3(n124), .S3(n111), .Z(n8814) );
  HS65_LL_IVX9 U13022 ( .A(n9135), .Z(n9127) );
  HS65_LL_IVX9 U13023 ( .A(n9134), .Z(n9128) );
  HS65_LL_NOR3AX2 U13024 ( .A(n8055), .B(n7765), .C(n8056), .Z(n8045) );
  HS65_LL_OAI21X3 U13025 ( .A(n343), .B(n7761), .C(n323), .Z(n8055) );
  HS65_LL_AOI12X2 U13026 ( .A(n399), .B(n368), .C(n8219), .Z(n8216) );
  HS65_LL_NOR2X6 U13027 ( .A(n630), .B(n627), .Z(n3691) );
  HS65_LL_NOR2X6 U13028 ( .A(n400), .B(n394), .Z(n8116) );
  HS65_LL_NOR2X6 U13029 ( .A(n327), .B(n329), .Z(n8356) );
  HS65_LL_NOR2X6 U13030 ( .A(n411), .B(n409), .Z(n3394) );
  HS65_LL_NAND4ABX3 U13031 ( .A(n8575), .B(n8576), .C(n8577), .D(n8578), .Z(
        n8560) );
  HS65_LL_NAND4ABX3 U13032 ( .A(n6743), .B(n6744), .C(n6745), .D(n6746), .Z(
        n6728) );
  HS65_LL_NAND4ABX3 U13033 ( .A(n5151), .B(n5152), .C(n5153), .D(n5154), .Z(
        n5136) );
  HS65_LL_NAND4ABX3 U13034 ( .A(n5383), .B(n5384), .C(n5385), .D(n5386), .Z(
        n5368) );
  HS65_LL_NAND4ABX3 U13035 ( .A(n6975), .B(n6976), .C(n6977), .D(n6978), .Z(
        n6960) );
  HS65_LL_NAND4ABX3 U13036 ( .A(n3636), .B(n3637), .C(n3638), .D(n3639), .Z(
        n3620) );
  HS65_LL_NOR2X6 U13037 ( .A(n275), .B(n274), .Z(n6544) );
  HS65_LL_NOR2X6 U13038 ( .A(n64), .B(n65), .Z(n6491) );
  HS65_LL_NOR2X6 U13039 ( .A(n233), .B(n232), .Z(n4898) );
  HS65_LL_NOR2X6 U13040 ( .A(n450), .B(n449), .Z(n4951) );
  HS65_LL_NOR2X6 U13041 ( .A(n502), .B(n501), .Z(n6416) );
  HS65_LL_NOR2X6 U13042 ( .A(n678), .B(n677), .Z(n4823) );
  HS65_LL_NAND2X7 U13043 ( .A(n158), .B(n179), .Z(n3029) );
  HS65_LL_NAND4ABX3 U13044 ( .A(n4818), .B(n5214), .C(n4859), .D(n5693), .Z(
        n5689) );
  HS65_LL_OAI21X3 U13045 ( .A(n696), .B(n691), .C(n666), .Z(n5693) );
  HS65_LL_NAND4ABX3 U13046 ( .A(n6411), .B(n6806), .C(n6452), .D(n7285), .Z(
        n7281) );
  HS65_LL_OAI21X3 U13047 ( .A(n520), .B(n515), .C(n490), .Z(n7285) );
  HS65_LL_NAND4ABX3 U13048 ( .A(n6642), .B(n6643), .C(n6644), .D(n6645), .Z(
        n6626) );
  HS65_LL_NAND4ABX3 U13049 ( .A(n5049), .B(n5050), .C(n5051), .D(n5052), .Z(
        n5033) );
  HS65_LL_NAND3AX6 U13050 ( .A(n3381), .B(n3382), .C(n3383), .Z(n3368) );
  HS65_LL_AOI12X2 U13051 ( .A(n420), .B(n3384), .C(n3385), .Z(n3383) );
  HS65_LL_NAND3AX6 U13052 ( .A(n3160), .B(n3161), .C(n3162), .Z(n3146) );
  HS65_LL_OAI21X3 U13053 ( .A(n661), .B(n3163), .C(n624), .Z(n3162) );
  HS65_LL_NAND3AX6 U13054 ( .A(n2960), .B(n2961), .C(n2962), .Z(n2945) );
  HS65_LL_OAI21X3 U13055 ( .A(n211), .B(n2963), .C(n201), .Z(n2962) );
  HS65_LL_NAND3X5 U13056 ( .A(n4713), .B(n4714), .C(n4715), .Z(n4697) );
  HS65_LL_AOI12X2 U13057 ( .A(n9), .B(n4716), .C(n4717), .Z(n4715) );
  HS65_LL_NAND3X5 U13058 ( .A(n6306), .B(n6307), .C(n6308), .Z(n6290) );
  HS65_LL_AOI12X2 U13059 ( .A(n531), .B(n6309), .C(n6310), .Z(n6308) );
  HS65_LL_CB4I6X9 U13060 ( .A(n567), .B(n568), .C(n531), .D(n6604), .Z(n6603)
         );
  HS65_LL_CB4I6X9 U13061 ( .A(n45), .B(n46), .C(n9), .D(n5011), .Z(n5010) );
  HS65_LL_CB4I6X9 U13062 ( .A(n524), .B(n525), .C(n489), .D(n6725), .Z(n6724)
         );
  HS65_LL_CB4I6X9 U13063 ( .A(n700), .B(n701), .C(n665), .D(n5133), .Z(n5132)
         );
  HS65_LL_CB4I6X9 U13064 ( .A(n88), .B(n91), .C(n69), .D(n6843), .Z(n6842) );
  HS65_LL_CB4I6X9 U13065 ( .A(n253), .B(n250), .C(n245), .D(n5251), .Z(n5250)
         );
  HS65_LL_CB4I6X9 U13066 ( .A(n470), .B(n467), .C(n462), .D(n5366), .Z(n5365)
         );
  HS65_LL_CB4I6X9 U13067 ( .A(n295), .B(n292), .C(n287), .D(n6958), .Z(n6957)
         );
  HS65_LL_BFX9 U13068 ( .A(n9148), .Z(n9146) );
  HS65_LL_BFX9 U13069 ( .A(n9148), .Z(n9147) );
  HS65_LL_MX41X7 U13070 ( .D0(n905), .S0(n889), .D1(n909), .S1(n890), .D2(n906), .S2(n884), .D3(n901), .S3(n885), .Z(n2550) );
  HS65_LL_MX41X7 U13071 ( .D0(n782), .S0(n766), .D1(n786), .S1(n767), .D2(n783), .S2(n761), .D3(n778), .S3(n762), .Z(n2174) );
  HS65_LL_MX41X7 U13072 ( .D0(n823), .S0(n807), .D1(n827), .S1(n808), .D2(n824), .S2(n802), .D3(n819), .S3(n803), .Z(n1798) );
  HS65_LL_MX41X7 U13073 ( .D0(n163), .S0(n143), .D1(n154), .S1(n175), .D2(n174), .S2(n151), .D3(n152), .S3(n167), .Z(n4097) );
  HS65_LL_MX41X7 U13074 ( .D0(n783), .S0(n761), .D1(n785), .S1(n768), .D2(n778), .S2(n771), .D3(n762), .S3(n792), .Z(n2008) );
  HS65_LL_MX41X7 U13075 ( .D0(n824), .S0(n802), .D1(n826), .S1(n809), .D2(n819), .S2(n812), .D3(n803), .S3(n833), .Z(n1632) );
  HS65_LL_MX41X7 U13076 ( .D0(n378), .S0(n383), .D1(n372), .S1(n396), .D2(n362), .S2(n399), .D3(n392), .S3(n377), .Z(n8200) );
  HS65_LL_MX41X7 U13077 ( .D0(n330), .S0(n344), .D1(n326), .S1(n356), .D2(n317), .S2(n350), .D3(n343), .S3(n329), .Z(n8503) );
  HS65_LL_MX41X7 U13078 ( .D0(n10), .S0(n29), .D1(n42), .S1(n25), .D2(n41), 
        .S2(n22), .D3(n23), .S3(n34), .Z(n5646) );
  HS65_LL_MX41X7 U13079 ( .D0(n532), .S0(n551), .D1(n564), .S1(n547), .D2(n563), .S2(n544), .D3(n545), .S3(n556), .Z(n7238) );
  HS65_LL_MX41X7 U13080 ( .D0(n258), .S0(n247), .D1(n264), .S1(n235), .D2(n267), .S2(n232), .D3(n263), .S3(n233), .Z(n5825) );
  HS65_LL_MX41X7 U13081 ( .D0(n475), .S0(n464), .D1(n481), .S1(n452), .D2(n484), .S2(n449), .D3(n480), .S3(n450), .Z(n5884) );
  HS65_LL_MX41X7 U13082 ( .D0(n684), .S0(n666), .D1(n697), .S1(n680), .D2(n696), .S2(n677), .D3(n689), .S3(n678), .Z(n5676) );
  HS65_LL_MX41X7 U13083 ( .D0(n73), .S0(n68), .D1(n78), .S1(n66), .D2(n81), 
        .S2(n65), .D3(n86), .S3(n64), .Z(n7417) );
  HS65_LL_MX41X7 U13084 ( .D0(n300), .S0(n289), .D1(n306), .S1(n277), .D2(n309), .S2(n274), .D3(n305), .S3(n275), .Z(n7476) );
  HS65_LL_MX41X7 U13085 ( .D0(n508), .S0(n490), .D1(n521), .S1(n504), .D2(n520), .S2(n501), .D3(n513), .S3(n502), .Z(n7268) );
  HS65_LL_MX41X7 U13086 ( .D0(n148), .S0(n174), .D1(n156), .S1(n178), .D2(n163), .S2(n149), .D3(n167), .S3(n155), .Z(n3547) );
  HS65_LL_MX41X7 U13087 ( .D0(n883), .S0(n907), .D1(n911), .S1(n895), .D2(n881), .S2(n902), .D3(n913), .S3(n2313), .Z(n2385) );
  HS65_LL_MX41X7 U13088 ( .D0(n193), .S0(n212), .D1(n201), .S1(n224), .D2(n218), .S2(n194), .D3(n213), .S3(n200), .Z(n3423) );
  HS65_LL_MX41X7 U13089 ( .D0(n320), .S0(n353), .D1(n343), .S1(n328), .D2(n329), .S2(n340), .D3(n327), .S3(n349), .Z(n8864) );
  HS65_LL_IVX9 U13090 ( .A(n7954), .Z(n321) );
  HS65_LL_OR3X9 U13091 ( .A(n1638), .B(n1639), .C(n1640), .Z(n1637) );
  HS65_LL_OR3X9 U13092 ( .A(n2390), .B(n2391), .C(n2392), .Z(n2389) );
  HS65_LL_OR3X9 U13093 ( .A(n1262), .B(n1263), .C(n1264), .Z(n1261) );
  HS65_LL_OR3X9 U13094 ( .A(n2014), .B(n2015), .C(n2016), .Z(n2013) );
  HS65_LL_OA12X9 U13095 ( .A(n7928), .B(n125), .C(n103), .Z(n7926) );
  HS65_LL_OA12X9 U13096 ( .A(n7830), .B(n605), .C(n583), .Z(n7828) );
  HS65_LL_OA12X9 U13097 ( .A(n4716), .B(n37), .C(n10), .Z(n5711) );
  HS65_LL_OA12X9 U13098 ( .A(n6309), .B(n559), .C(n532), .Z(n7303) );
  HS65_LL_CBI4I6X5 U13099 ( .A(n888), .B(n2428), .C(n908), .D(n2523), .Z(n2503) );
  HS65_LL_OA12X9 U13100 ( .A(n2346), .B(n913), .C(n892), .Z(n2523) );
  HS65_LL_OA12X9 U13101 ( .A(n3236), .B(n152), .C(n174), .Z(n3911) );
  HS65_LL_AO12X9 U13102 ( .A(n405), .B(n443), .C(n3169), .Z(n3168) );
  HS65_LL_AO12X9 U13103 ( .A(n201), .B(n218), .C(n2942), .Z(n2941) );
  HS65_LL_AO12X9 U13104 ( .A(n624), .B(n652), .C(n3143), .Z(n3142) );
  HS65_LL_AO12X9 U13105 ( .A(n156), .B(n163), .C(n3018), .Z(n3017) );
  HS65_LL_AO12X9 U13106 ( .A(n19), .B(n29), .C(n4542), .Z(n4541) );
  HS65_LL_AO12X9 U13107 ( .A(n541), .B(n551), .C(n6135), .Z(n6134) );
  HS65_LL_AO12X9 U13108 ( .A(n236), .B(n258), .C(n4740), .Z(n4739) );
  HS65_LL_AO12X9 U13109 ( .A(n453), .B(n475), .C(n4766), .Z(n4765) );
  HS65_LL_AO12X9 U13110 ( .A(n278), .B(n300), .C(n6359), .Z(n6358) );
  HS65_LL_AO12X9 U13111 ( .A(n59), .B(n73), .C(n6320), .Z(n6319) );
  HS65_LL_AO12X9 U13112 ( .A(n498), .B(n508), .C(n6212), .Z(n6211) );
  HS65_LL_AO12X9 U13113 ( .A(n674), .B(n684), .C(n4619), .Z(n4618) );
  HS65_LL_OA12X9 U13114 ( .A(n3101), .B(n215), .C(n189), .Z(n4180) );
  HS65_LL_OA12X9 U13115 ( .A(n8110), .B(n399), .C(n363), .Z(n8969) );
  HS65_LL_OA12X9 U13116 ( .A(n4980), .B(n478), .C(n464), .Z(n5624) );
  HS65_LL_OA12X9 U13117 ( .A(n4927), .B(n261), .C(n247), .Z(n5599) );
  HS65_LL_OA12X9 U13118 ( .A(n6573), .B(n303), .C(n289), .Z(n7216) );
  HS65_LL_OA12X9 U13119 ( .A(n4854), .B(n692), .C(n666), .Z(n5773) );
  HS65_LL_OA12X9 U13120 ( .A(n6447), .B(n516), .C(n490), .Z(n7365) );
  HS65_LL_OA12X9 U13121 ( .A(n6520), .B(n85), .C(n68), .Z(n7191) );
  HS65_LL_OA12X9 U13122 ( .A(n8343), .B(n350), .C(n320), .Z(n8909) );
  HS65_LL_OA12X9 U13123 ( .A(n3257), .B(n170), .C(n143), .Z(n4118) );
  HS65_LL_AO12X9 U13124 ( .A(n373), .B(n395), .C(n7973), .Z(n7972) );
  HS65_LL_AO12X9 U13125 ( .A(n323), .B(n353), .C(n8041), .Z(n8040) );
  HS65_LL_OA12X9 U13126 ( .A(n3384), .B(n437), .C(n422), .Z(n4032) );
  HS65_LL_OA12X9 U13127 ( .A(n3330), .B(n654), .C(n640), .Z(n4009) );
  HS65_LL_OA12X9 U13128 ( .A(n7864), .B(n371), .C(n397), .Z(n7863) );
  HS65_LL_OA12X9 U13129 ( .A(n6120), .B(n497), .C(n515), .Z(n6119) );
  HS65_LL_OA12X9 U13130 ( .A(n4527), .B(n673), .C(n691), .Z(n4526) );
  HS65_LL_OA12X9 U13131 ( .A(n4458), .B(n237), .C(n262), .Z(n4592) );
  HS65_LL_OA12X9 U13132 ( .A(n6090), .B(n279), .C(n304), .Z(n6202) );
  HS65_LL_OA12X9 U13133 ( .A(n6051), .B(n58), .C(n84), .Z(n6185) );
  HS65_LL_OA12X9 U13134 ( .A(n4497), .B(n454), .C(n479), .Z(n4609) );
  HS65_LL_OA12X9 U13135 ( .A(n1114), .B(n871), .C(n845), .Z(n1142) );
  HS65_LL_OA12X9 U13136 ( .A(n1866), .B(n789), .C(n763), .Z(n1894) );
  HS65_LL_OA12X9 U13137 ( .A(n2242), .B(n912), .C(n886), .Z(n2270) );
  HS65_LL_OA12X9 U13138 ( .A(n1490), .B(n830), .C(n804), .Z(n1518) );
  HS65_LL_OA12X9 U13139 ( .A(n2834), .B(n407), .C(n438), .Z(n2991) );
  HS65_LL_OA12X9 U13140 ( .A(n2912), .B(n155), .C(n168), .Z(n2911) );
  HS65_LL_OA12X9 U13141 ( .A(n2886), .B(n626), .C(n655), .Z(n2980) );
  HS65_LL_OA12X9 U13142 ( .A(n2869), .B(n200), .C(n214), .Z(n2868) );
  HS65_LL_OA12X9 U13143 ( .A(n7946), .B(n324), .C(n352), .Z(n7945) );
  HS65_LL_OA12X9 U13144 ( .A(n7833), .B(n591), .C(n606), .Z(n8006) );
  HS65_LL_OA12X9 U13145 ( .A(n7872), .B(n111), .C(n126), .Z(n8019) );
  HS65_LL_OA12X9 U13146 ( .A(n6080), .B(n540), .C(n558), .Z(n6079) );
  HS65_LL_OA12X9 U13147 ( .A(n4487), .B(n18), .C(n36), .Z(n4486) );
  HS65_LL_IVX9 U13148 ( .A(n6149), .Z(n534) );
  HS65_LL_IVX9 U13149 ( .A(n4556), .Z(n12) );
  HS65_LL_OA12X9 U13150 ( .A(n349), .B(n8619), .C(n324), .Z(n8617) );
  HS65_LL_OA12X9 U13151 ( .A(n398), .B(n8492), .C(n371), .Z(n8659) );
  HS65_LL_IVX9 U13152 ( .A(n8717), .Z(n589) );
  HS65_LL_AND3X9 U13153 ( .A(n5141), .B(n4634), .C(n5159), .Z(n5686) );
  HS65_LL_AND3X9 U13154 ( .A(n6733), .B(n6227), .C(n6751), .Z(n7278) );
  HS65_LL_BFX9 U13155 ( .A(n9133), .Z(n9132) );
  HS65_LL_NAND4X9 U13156 ( .A(n5080), .B(n5081), .C(n5082), .D(n5083), .Z(
        n5074) );
  HS65_LL_NAND4X9 U13157 ( .A(n6673), .B(n6674), .C(n6675), .D(n6676), .Z(
        n6667) );
  HS65_LL_NAND2X7 U13158 ( .A(n2582), .B(n2583), .Z(n2246) );
  HS65_LL_NAND2X7 U13159 ( .A(n1830), .B(n1831), .Z(n1494) );
  HS65_LL_NAND2X7 U13160 ( .A(n1454), .B(n1455), .Z(n1118) );
  HS65_LL_NAND2X7 U13161 ( .A(n2206), .B(n2207), .Z(n1870) );
  HS65_LL_NAND2X7 U13162 ( .A(n4270), .B(n4271), .Z(n2882) );
  HS65_LL_NAND2X7 U13163 ( .A(n8988), .B(n8989), .Z(n7851) );
  HS65_LL_NAND2X7 U13164 ( .A(n4137), .B(n4152), .Z(n2918) );
  HS65_LL_NAND2X7 U13165 ( .A(n4212), .B(n4202), .Z(n2860) );
  HS65_LL_NOR4ABX2 U13166 ( .A(n7994), .B(n7995), .C(n7996), .D(n7997), .Z(
        n2780) );
  HS65_LL_CBI4I1X5 U13167 ( .A(n7686), .B(n7806), .C(n7618), .D(n8003), .Z(
        n7996) );
  HS65_LL_CBI4I6X5 U13168 ( .A(n585), .B(n7699), .C(n616), .D(n8004), .Z(n7995) );
  HS65_LL_AOI212X4 U13169 ( .A(n600), .B(n580), .C(n587), .D(n610), .E(n8006), 
        .Z(n7994) );
  HS65_LL_NOR4ABX2 U13170 ( .A(n3886), .B(n3887), .C(n3888), .D(n3889), .Z(
        n2666) );
  HS65_LL_CBI4I1X5 U13171 ( .A(n2933), .B(n3095), .C(n2856), .D(n3514), .Z(
        n3888) );
  HS65_LL_CBI4I1X5 U13172 ( .A(n3890), .B(n3097), .C(n2859), .D(n3891), .Z(
        n3889) );
  HS65_LL_AOI212X4 U13173 ( .A(n215), .B(n200), .C(n201), .D(n3897), .E(n3898), 
        .Z(n3886) );
  HS65_LL_NOR4ABX2 U13174 ( .A(n8007), .B(n8008), .C(n8009), .D(n8010), .Z(
        n2804) );
  HS65_LL_CBI4I1X5 U13175 ( .A(n7724), .B(n7869), .C(n7659), .D(n8016), .Z(
        n8009) );
  HS65_LL_CBI4I6X5 U13176 ( .A(n105), .B(n7737), .C(n136), .D(n8017), .Z(n8008) );
  HS65_LL_AOI212X4 U13177 ( .A(n120), .B(n100), .C(n107), .D(n130), .E(n8019), 
        .Z(n8007) );
  HS65_LL_NOR4ABX2 U13178 ( .A(n7865), .B(n7866), .C(n7867), .D(n7868), .Z(
        n2805) );
  HS65_LL_NAND4ABX3 U13179 ( .A(n7876), .B(n7877), .C(n7878), .D(n7879), .Z(
        n7867) );
  HS65_LL_OAI212X5 U13180 ( .A(n7714), .B(n7869), .C(n7650), .D(n7870), .E(
        n7871), .Z(n7868) );
  HS65_LL_AOI212X4 U13181 ( .A(n105), .B(n126), .C(n119), .D(n113), .E(n7881), 
        .Z(n7866) );
  HS65_LL_NOR4ABX2 U13182 ( .A(n4655), .B(n4656), .C(n4657), .D(n4658), .Z(
        n2770) );
  HS65_LL_NAND4ABX3 U13183 ( .A(n4663), .B(n4664), .C(n4665), .D(n4666), .Z(
        n4657) );
  HS65_LL_OAI212X5 U13184 ( .A(n4659), .B(n4550), .C(n4660), .D(n4661), .E(
        n4662), .Z(n4658) );
  HS65_LL_AOI212X4 U13185 ( .A(n19), .B(n38), .C(n47), .D(n22), .E(n4669), .Z(
        n4656) );
  HS65_LL_NOR4ABX2 U13186 ( .A(n6248), .B(n6249), .C(n6250), .D(n6251), .Z(
        n2762) );
  HS65_LL_NAND4ABX3 U13187 ( .A(n6256), .B(n6257), .C(n6258), .D(n6259), .Z(
        n6250) );
  HS65_LL_OAI212X5 U13188 ( .A(n6252), .B(n6143), .C(n6253), .D(n6254), .E(
        n6255), .Z(n6251) );
  HS65_LL_AOI212X4 U13189 ( .A(n541), .B(n560), .C(n569), .D(n544), .E(n6262), 
        .Z(n6249) );
  HS65_LL_NOR4ABX2 U13190 ( .A(n3287), .B(n3288), .C(n3289), .D(n3290), .Z(
        n2641) );
  HS65_LL_OAI212X5 U13191 ( .A(n3291), .B(n2884), .C(n3292), .D(n3293), .E(
        n3294), .Z(n3290) );
  HS65_LL_NAND4ABX3 U13192 ( .A(n3295), .B(n3296), .C(n3297), .D(n3298), .Z(
        n3289) );
  HS65_LL_AOI212X4 U13193 ( .A(n624), .B(n657), .C(n645), .D(n628), .E(n3300), 
        .Z(n3288) );
  HS65_LL_IVX9 U13194 ( .A(n8039), .Z(n351) );
  HS65_LL_NOR4ABX2 U13195 ( .A(n6187), .B(n6188), .C(n6189), .D(n6190), .Z(
        n2812) );
  HS65_LL_CBI4I6X5 U13196 ( .A(n276), .B(n6199), .C(n301), .D(n6200), .Z(n6188) );
  HS65_LL_CBI4I1X5 U13197 ( .A(n6196), .B(n6086), .C(n6197), .D(n6198), .Z(
        n6189) );
  HS65_LL_AOI212X4 U13198 ( .A(n295), .B(n285), .C(n309), .D(n277), .E(n6202), 
        .Z(n6187) );
  HS65_LL_NOR4ABX2 U13199 ( .A(n4594), .B(n4595), .C(n4596), .D(n4597), .Z(
        n2820) );
  HS65_LL_CBI4I6X5 U13200 ( .A(n451), .B(n4606), .C(n476), .D(n4607), .Z(n4595) );
  HS65_LL_CBI4I1X5 U13201 ( .A(n4603), .B(n4493), .C(n4604), .D(n4605), .Z(
        n4596) );
  HS65_LL_AOI212X4 U13202 ( .A(n470), .B(n460), .C(n484), .D(n452), .E(n4609), 
        .Z(n4594) );
  HS65_LL_NOR4ABX2 U13203 ( .A(n6061), .B(n6062), .C(n6063), .D(n6064), .Z(
        n2764) );
  HS65_LL_CBI4I6X5 U13204 ( .A(n546), .B(n6074), .C(n552), .D(n6075), .Z(n6062) );
  HS65_LL_CBI4I1X5 U13205 ( .A(n6070), .B(n6071), .C(n6072), .D(n6073), .Z(
        n6063) );
  HS65_LL_AOI212X4 U13206 ( .A(n539), .B(n567), .C(n563), .D(n547), .E(n6079), 
        .Z(n6061) );
  HS65_LL_NOR4ABX2 U13207 ( .A(n4468), .B(n4469), .C(n4470), .D(n4471), .Z(
        n2772) );
  HS65_LL_CBI4I6X5 U13208 ( .A(n24), .B(n4481), .C(n30), .D(n4482), .Z(n4469)
         );
  HS65_LL_CBI4I1X5 U13209 ( .A(n4477), .B(n4478), .C(n4479), .D(n4480), .Z(
        n4470) );
  HS65_LL_AOI212X4 U13210 ( .A(n17), .B(n45), .C(n41), .D(n25), .E(n4486), .Z(
        n4468) );
  HS65_LL_NOR4ABX2 U13211 ( .A(n7842), .B(n7843), .C(n7844), .D(n7845), .Z(
        n2756) );
  HS65_LL_CBI4I1X5 U13212 ( .A(n7846), .B(n7847), .C(n7848), .D(n7849), .Z(
        n7845) );
  HS65_LL_CBI4I1X5 U13213 ( .A(n7850), .B(n7851), .C(n7852), .D(n7853), .Z(
        n7844) );
  HS65_LL_AOI212X4 U13214 ( .A(n384), .B(n370), .C(n376), .D(n389), .E(n7863), 
        .Z(n7842) );
  HS65_LL_NOR4ABX2 U13215 ( .A(n6463), .B(n6464), .C(n6465), .D(n6466), .Z(
        n2786) );
  HS65_LL_NAND4ABX3 U13216 ( .A(n6471), .B(n6472), .C(n6473), .D(n6474), .Z(
        n6465) );
  HS65_LL_OAI212X5 U13217 ( .A(n6467), .B(n6048), .C(n6468), .D(n6469), .E(
        n6470), .Z(n6466) );
  HS65_LL_AOI212X4 U13218 ( .A(n59), .B(n80), .C(n89), .D(n65), .E(n6477), .Z(
        n6464) );
  HS65_LL_NOR4ABX2 U13219 ( .A(n4870), .B(n4871), .C(n4872), .D(n4873), .Z(
        n2794) );
  HS65_LL_NAND4ABX3 U13220 ( .A(n4878), .B(n4879), .C(n4880), .D(n4881), .Z(
        n4872) );
  HS65_LL_OAI212X5 U13221 ( .A(n4874), .B(n4455), .C(n4875), .D(n4876), .E(
        n4877), .Z(n4873) );
  HS65_LL_AOI212X4 U13222 ( .A(n236), .B(n266), .C(n252), .D(n232), .E(n4884), 
        .Z(n4871) );
  HS65_LL_NOR4ABX2 U13223 ( .A(n8873), .B(n8874), .C(n8875), .D(n8876), .Z(
        n2620) );
  HS65_LL_CBI4I1X5 U13224 ( .A(n7953), .B(n7942), .C(n7768), .D(n8877), .Z(
        n8876) );
  HS65_LL_CBI4I1X5 U13225 ( .A(n7940), .B(n8630), .C(n8034), .D(n8578), .Z(
        n8875) );
  HS65_LL_AOI222X2 U13226 ( .A(n332), .B(n349), .C(n323), .D(n8933), .E(n353), 
        .F(n327), .Z(n8873) );
  HS65_LL_NOR4ABX2 U13227 ( .A(n3931), .B(n3932), .C(n3933), .D(n3934), .Z(
        n2659) );
  HS65_LL_CBI4I1X5 U13228 ( .A(n3135), .B(n2883), .C(n2969), .D(n3753), .Z(
        n3933) );
  HS65_LL_CBI4I1X5 U13229 ( .A(n3935), .B(n2881), .C(n2972), .D(n3936), .Z(
        n3934) );
  HS65_LL_AOI212X4 U13230 ( .A(n654), .B(n626), .C(n624), .D(n2895), .E(n3951), 
        .Z(n3931) );
  HS65_LL_NOR4ABX2 U13231 ( .A(n2851), .B(n2852), .C(n2853), .D(n2854), .Z(
        n2637) );
  HS65_LL_CBI4I1X5 U13232 ( .A(n2859), .B(n2860), .C(n2861), .D(n2862), .Z(
        n2853) );
  HS65_LL_CBI4I1X5 U13233 ( .A(n2855), .B(n2856), .C(n2857), .D(n2858), .Z(
        n2854) );
  HS65_LL_AOI212X4 U13234 ( .A(n194), .B(n224), .C(n199), .D(n212), .E(n2868), 
        .Z(n2851) );
  HS65_LL_NOR4ABX2 U13235 ( .A(n2964), .B(n2965), .C(n2966), .D(n2967), .Z(
        n2627) );
  HS65_LL_CBI4I1X5 U13236 ( .A(n2968), .B(n2969), .C(n2970), .D(n2971), .Z(
        n2967) );
  HS65_LL_CBI4I1X5 U13237 ( .A(n2972), .B(n2882), .C(n2973), .D(n2974), .Z(
        n2966) );
  HS65_LL_AOI212X4 U13238 ( .A(n635), .B(n646), .C(n630), .D(n659), .E(n2980), 
        .Z(n2964) );
  HS65_LL_NOR4ABX2 U13239 ( .A(n7089), .B(n7090), .C(n7091), .D(n7092), .Z(
        n2759) );
  HS65_LL_CB4I6X9 U13240 ( .A(n555), .B(n553), .C(n540), .D(n6642), .Z(n7091)
         );
  HS65_LL_CBI4I1X5 U13241 ( .A(n6072), .B(n7093), .C(n7094), .D(n7095), .Z(
        n7092) );
  HS65_LL_AOI222X2 U13242 ( .A(n537), .B(n556), .C(n541), .D(n7108), .E(n545), 
        .F(n551), .Z(n7089) );
  HS65_LL_NOR4ABX2 U13243 ( .A(n5497), .B(n5498), .C(n5499), .D(n5500), .Z(
        n2767) );
  HS65_LL_CB4I6X9 U13244 ( .A(n33), .B(n31), .C(n18), .D(n5049), .Z(n5499) );
  HS65_LL_CBI4I1X5 U13245 ( .A(n4479), .B(n5501), .C(n5502), .D(n5503), .Z(
        n5500) );
  HS65_LL_AOI222X2 U13246 ( .A(n15), .B(n34), .C(n19), .D(n5516), .E(n23), .F(
        n29), .Z(n5497) );
  HS65_LL_NOR4ABX2 U13247 ( .A(n3996), .B(n3997), .C(n3998), .D(n3999), .Z(
        n2663) );
  HS65_LL_CB4I6X9 U13248 ( .A(n650), .B(n649), .C(n626), .D(n3746), .Z(n3998)
         );
  HS65_LL_CBI4I1X5 U13249 ( .A(n2973), .B(n3140), .C(n3342), .D(n4000), .Z(
        n3999) );
  HS65_LL_AOI222X2 U13250 ( .A(n636), .B(n656), .C(n624), .D(n4019), .E(n629), 
        .F(n652), .Z(n3996) );
  HS65_LL_IVX9 U13251 ( .A(n8049), .Z(n348) );
  HS65_LL_NOR4ABX2 U13252 ( .A(n7230), .B(n7231), .C(n7232), .D(n7233), .Z(
        n2758) );
  HS65_LL_MX41X7 U13253 ( .D0(n559), .S0(n538), .D1(n569), .S1(n544), .D2(n545), .S2(n558), .D3(n539), .S3(n6154), .Z(n7233) );
  HS65_LL_MX41X7 U13254 ( .D0(n557), .S0(n6074), .D1(n531), .S1(n553), .D2(
        n536), .S2(n568), .D3(n555), .S3(n541), .Z(n7232) );
  HS65_LL_NOR4ABX2 U13255 ( .A(n6631), .B(n6611), .C(n7234), .D(n6147), .Z(
        n7231) );
  HS65_LL_IVX9 U13256 ( .A(n7981), .Z(n387) );
  HS65_LL_NAND4ABX3 U13257 ( .A(n7666), .B(n7667), .C(n7668), .D(n7669), .Z(
        n2774) );
  HS65_LL_MX41X7 U13258 ( .D0(n605), .S0(n576), .D1(n588), .S1(n602), .D2(n586), .S2(n606), .D3(n580), .S3(n7700), .Z(n7667) );
  HS65_LL_MX41X7 U13259 ( .D0(n607), .S0(n7699), .D1(n584), .S1(n617), .D2(
        n579), .S2(n603), .D3(n614), .S3(n592), .Z(n7666) );
  HS65_LL_NOR4ABX2 U13260 ( .A(n7670), .B(n7671), .C(n7672), .D(n7673), .Z(
        n7669) );
  HS65_LL_NAND4ABX3 U13261 ( .A(n8631), .B(n8632), .C(n8633), .D(n8634), .Z(
        n2757) );
  HS65_LL_OAI212X5 U13262 ( .A(n7851), .B(n7751), .C(n8106), .D(n7861), .E(
        n8657), .Z(n8632) );
  HS65_LL_NAND4ABX3 U13263 ( .A(n8659), .B(n8298), .C(n8262), .D(n8660), .Z(
        n8631) );
  HS65_LL_AOI212X4 U13264 ( .A(n378), .B(n397), .C(n372), .D(n386), .E(n8635), 
        .Z(n8634) );
  HS65_LL_NAND4ABX3 U13265 ( .A(n2870), .B(n2871), .C(n2872), .D(n2873), .Z(
        n2630) );
  HS65_LL_NAND4ABX3 U13266 ( .A(n2891), .B(n2892), .C(n2893), .D(n2894), .Z(
        n2870) );
  HS65_LL_OAI212X5 U13267 ( .A(n2881), .B(n2882), .C(n2883), .D(n2884), .E(
        n2885), .Z(n2871) );
  HS65_LL_AOI212X4 U13268 ( .A(n631), .B(n655), .C(n625), .D(n648), .E(n2874), 
        .Z(n2873) );
  HS65_LL_NAND4ABX3 U13269 ( .A(n5757), .B(n5758), .C(n5759), .D(n5760), .Z(
        n3533) );
  HS65_LL_OAI212X5 U13270 ( .A(n4850), .B(n4534), .C(n4626), .D(n4848), .E(
        n5815), .Z(n5758) );
  HS65_LL_NAND4ABX3 U13271 ( .A(n5170), .B(n5218), .C(n5817), .D(n5818), .Z(
        n5757) );
  HS65_LL_AOI212X4 U13272 ( .A(n679), .B(n691), .C(n675), .D(n699), .E(n5761), 
        .Z(n5760) );
  HS65_LL_NAND4ABX3 U13273 ( .A(n7349), .B(n7350), .C(n7351), .D(n7352), .Z(
        n3208) );
  HS65_LL_OAI212X5 U13274 ( .A(n6443), .B(n6127), .C(n6219), .D(n6441), .E(
        n7407), .Z(n7350) );
  HS65_LL_NAND4ABX3 U13275 ( .A(n6762), .B(n6810), .C(n7409), .D(n7410), .Z(
        n7349) );
  HS65_LL_AOI212X4 U13276 ( .A(n503), .B(n515), .C(n499), .D(n523), .E(n7353), 
        .Z(n7352) );
  HS65_LL_NOR4ABX2 U13277 ( .A(n7411), .B(n7412), .C(n7413), .D(n7414), .Z(
        n2782) );
  HS65_LL_MX41X7 U13278 ( .D0(n85), .S0(n54), .D1(n89), .S1(n65), .D2(n64), 
        .S2(n84), .D3(n56), .S3(n6338), .Z(n7414) );
  HS65_LL_MX41X7 U13279 ( .D0(n83), .S0(n6182), .D1(n69), .S1(n74), .D2(n57), 
        .S2(n91), .D3(n76), .S3(n59), .Z(n7413) );
  HS65_LL_NOR4ABX2 U13280 ( .A(n6869), .B(n7415), .C(n6851), .D(n6331), .Z(
        n7412) );
  HS65_LL_NOR4ABX2 U13281 ( .A(n8611), .B(n8612), .C(n8613), .D(n8614), .Z(
        n3005) );
  HS65_LL_OAI212X5 U13282 ( .A(n7952), .B(n7769), .C(n8339), .D(n7943), .E(
        n8615), .Z(n8614) );
  HS65_LL_NAND4ABX3 U13283 ( .A(n8617), .B(n8523), .C(n8564), .D(n8618), .Z(
        n8613) );
  HS65_LL_AOI212X4 U13284 ( .A(n330), .B(n352), .C(n326), .D(n347), .E(n8620), 
        .Z(n8612) );
  HS65_LL_IVX9 U13285 ( .A(n7846), .Z(n362) );
  HS65_LL_NAND4ABX3 U13286 ( .A(n7778), .B(n7779), .C(n7780), .D(n7781), .Z(
        n2781) );
  HS65_LL_NAND4ABX3 U13287 ( .A(n7837), .B(n7838), .C(n7839), .D(n7840), .Z(
        n7778) );
  HS65_LL_OAI212X5 U13288 ( .A(n7676), .B(n7806), .C(n7630), .D(n7831), .E(
        n7832), .Z(n7779) );
  HS65_LL_AOI212X4 U13289 ( .A(n585), .B(n606), .C(n599), .D(n593), .E(n7782), 
        .Z(n7781) );
  HS65_LL_NOR4ABX2 U13290 ( .A(n7065), .B(n7096), .C(n7097), .D(n7098), .Z(
        n7090) );
  HS65_LL_OAI212X5 U13291 ( .A(n7099), .B(n6143), .C(n7100), .D(n6078), .E(
        n7101), .Z(n7098) );
  HS65_LL_NOR4ABX2 U13292 ( .A(n5473), .B(n5504), .C(n5505), .D(n5506), .Z(
        n5498) );
  HS65_LL_OAI212X5 U13293 ( .A(n5507), .B(n4550), .C(n5508), .D(n4485), .E(
        n5509), .Z(n5506) );
  HS65_LL_NAND4ABX3 U13294 ( .A(n5695), .B(n5696), .C(n5697), .D(n5698), .Z(
        n2773) );
  HS65_LL_OAI212X5 U13295 ( .A(n4478), .B(n4712), .C(n4709), .D(n4550), .E(
        n5753), .Z(n5696) );
  HS65_LL_NAND4ABX3 U13296 ( .A(n5048), .B(n5112), .C(n5755), .D(n5756), .Z(
        n5695) );
  HS65_LL_AOI212X4 U13297 ( .A(n24), .B(n36), .C(n44), .D(n20), .E(n5699), .Z(
        n5698) );
  HS65_LL_NAND4ABX3 U13298 ( .A(n7287), .B(n7288), .C(n7289), .D(n7290), .Z(
        n2765) );
  HS65_LL_OAI212X5 U13299 ( .A(n6071), .B(n6305), .C(n6302), .D(n6143), .E(
        n7345), .Z(n7288) );
  HS65_LL_NAND4ABX3 U13300 ( .A(n6641), .B(n6705), .C(n7347), .D(n7348), .Z(
        n7287) );
  HS65_LL_AOI212X4 U13301 ( .A(n546), .B(n558), .C(n566), .D(n542), .E(n7291), 
        .Z(n7290) );
  HS65_LL_NAND4ABX3 U13302 ( .A(n7203), .B(n7204), .C(n7205), .D(n7206), .Z(
        n2807) );
  HS65_LL_CB4I6X9 U13303 ( .A(n299), .B(n298), .C(n279), .D(n6994), .Z(n7203)
         );
  HS65_LL_AOI222X2 U13304 ( .A(n305), .B(n286), .C(n278), .D(n7228), .E(n300), 
        .F(n275), .Z(n7205) );
  HS65_LL_CBI4I1X5 U13305 ( .A(n6197), .B(n7146), .C(n7222), .D(n7229), .Z(
        n7204) );
  HS65_LL_NAND4ABX3 U13306 ( .A(n4102), .B(n4103), .C(n4104), .D(n4105), .Z(
        n2682) );
  HS65_LL_OAI212X5 U13307 ( .A(n3253), .B(n2918), .C(n3032), .D(n3251), .E(
        n4160), .Z(n4103) );
  HS65_LL_NAND4ABX3 U13308 ( .A(n3635), .B(n3567), .C(n4162), .D(n4163), .Z(
        n4102) );
  HS65_LL_AOI212X4 U13309 ( .A(n168), .B(n153), .C(n158), .D(n177), .E(n4106), 
        .Z(n4105) );
  HS65_LL_IVX9 U13310 ( .A(n1180), .Z(n843) );
  HS65_LL_IVX9 U13311 ( .A(n1932), .Z(n761) );
  HS65_LL_IVX9 U13312 ( .A(n2308), .Z(n884) );
  HS65_LL_IVX9 U13313 ( .A(n1556), .Z(n802) );
  HS65_LL_IVX9 U13314 ( .A(n2958), .Z(n225) );
  HS65_LL_IVX9 U13315 ( .A(n3185), .Z(n431) );
  HS65_LL_OAI212X5 U13316 ( .A(n1407), .B(n1116), .C(n1317), .D(n1143), .E(
        n1408), .Z(n1406) );
  HS65_LL_OAI21X3 U13317 ( .A(n866), .B(n873), .C(n855), .Z(n1408) );
  HS65_LL_NOR3X4 U13318 ( .A(n841), .B(n850), .C(n843), .Z(n1407) );
  HS65_LL_OAI212X5 U13319 ( .A(n2159), .B(n1868), .C(n2069), .D(n1895), .E(
        n2160), .Z(n2158) );
  HS65_LL_OAI21X3 U13320 ( .A(n784), .B(n791), .C(n773), .Z(n2160) );
  HS65_LL_NOR3X4 U13321 ( .A(n759), .B(n768), .C(n761), .Z(n2159) );
  HS65_LL_OAI212X5 U13322 ( .A(n1783), .B(n1492), .C(n1693), .D(n1519), .E(
        n1784), .Z(n1782) );
  HS65_LL_NOR3X4 U13323 ( .A(n800), .B(n809), .C(n802), .Z(n1783) );
  HS65_LL_OAI21X3 U13324 ( .A(n825), .B(n832), .C(n814), .Z(n1784) );
  HS65_LL_IVX9 U13325 ( .A(n3158), .Z(n644) );
  HS65_LL_NAND4ABX3 U13326 ( .A(n5638), .B(n5639), .C(n5640), .D(n5641), .Z(
        n2766) );
  HS65_LL_NOR4ABX2 U13327 ( .A(n5038), .B(n5018), .C(n5642), .D(n4554), .Z(
        n5641) );
  HS65_LL_MX41X7 U13328 ( .D0(n35), .S0(n4481), .D1(n9), .S1(n31), .D2(n14), 
        .S2(n46), .D3(n33), .S3(n19), .Z(n5638) );
  HS65_LL_MX41X7 U13329 ( .D0(n37), .S0(n16), .D1(n47), .S1(n22), .D2(n23), 
        .S2(n36), .D3(n17), .S3(n4561), .Z(n5639) );
  HS65_LL_NAND4ABX3 U13330 ( .A(n8995), .B(n8996), .C(n8997), .D(n8998), .Z(
        n2776) );
  HS65_LL_CBI4I1X5 U13331 ( .A(n7622), .B(n7831), .C(n8397), .D(n8700), .Z(
        n8995) );
  HS65_LL_AOI212X4 U13332 ( .A(n591), .B(n605), .C(n592), .D(n7841), .E(n9050), 
        .Z(n8997) );
  HS65_LL_CBI4I1X5 U13333 ( .A(n8719), .B(n7676), .C(n7686), .D(n9052), .Z(
        n8996) );
  HS65_LL_NAND4ABX3 U13334 ( .A(n4164), .B(n4165), .C(n4166), .D(n4167), .Z(
        n2722) );
  HS65_LL_NAND4ABX3 U13335 ( .A(n3503), .B(n3446), .C(n4224), .D(n4225), .Z(
        n4164) );
  HS65_LL_OAI212X5 U13336 ( .A(n3097), .B(n2860), .C(n3095), .D(n2956), .E(
        n4222), .Z(n4165) );
  HS65_LL_AOI212X4 U13337 ( .A(n198), .B(n214), .C(n203), .D(n223), .E(n4168), 
        .Z(n4167) );
  HS65_LL_NAND4ABX3 U13338 ( .A(n5819), .B(n5820), .C(n5821), .D(n5822), .Z(
        n2790) );
  HS65_LL_NOR4ABX2 U13339 ( .A(n5277), .B(n5823), .C(n5259), .D(n4750), .Z(
        n5822) );
  HS65_LL_MX41X7 U13340 ( .D0(n260), .S0(n4589), .D1(n245), .S1(n256), .D2(
        n241), .S2(n250), .D3(n257), .S3(n236), .Z(n5819) );
  HS65_LL_MX41X7 U13341 ( .D0(n261), .S0(n242), .D1(n252), .S1(n232), .D2(n233), .S2(n262), .D3(n243), .S3(n4757), .Z(n5820) );
  HS65_LL_NAND4ABX3 U13342 ( .A(n7642), .B(n7643), .C(n7644), .D(n7645), .Z(
        n2799) );
  HS65_LL_CBI4I1X5 U13343 ( .A(n7662), .B(n7663), .C(n7664), .D(n7665), .Z(
        n7642) );
  HS65_LL_CBI4I1X5 U13344 ( .A(n7659), .B(n7656), .C(n7660), .D(n7661), .Z(
        n7643) );
  HS65_LL_AOI222X2 U13345 ( .A(n124), .B(n98), .C(n112), .D(n7655), .E(n135), 
        .F(n106), .Z(n7644) );
  HS65_LL_NAND4ABX3 U13346 ( .A(n7156), .B(n7157), .C(n7158), .D(n7159), .Z(
        n3007) );
  HS65_LL_CB4I6X9 U13347 ( .A(n512), .B(n510), .C(n497), .D(n6763), .Z(n7156)
         );
  HS65_LL_AOI222X2 U13348 ( .A(n513), .B(n494), .C(n498), .D(n7174), .E(n508), 
        .F(n502), .Z(n7158) );
  HS65_LL_CBI4I1X5 U13349 ( .A(n6128), .B(n7171), .C(n7173), .D(n7175), .Z(
        n7157) );
  HS65_LL_IVX9 U13350 ( .A(n1861), .Z(n765) );
  HS65_LL_NOR4ABX2 U13351 ( .A(n8849), .B(n8855), .C(n8623), .D(n8878), .Z(
        n8874) );
  HS65_LL_OAI212X5 U13352 ( .A(n8039), .B(n7943), .C(n8540), .D(n8527), .E(
        n7772), .Z(n8878) );
  HS65_LL_IVX9 U13353 ( .A(n1109), .Z(n847) );
  HS65_LL_IVX9 U13354 ( .A(n2237), .Z(n888) );
  HS65_LL_IVX9 U13355 ( .A(n1485), .Z(n806) );
  HS65_LL_NAND4ABX3 U13356 ( .A(n5564), .B(n5565), .C(n5566), .D(n5567), .Z(
        n3210) );
  HS65_LL_CB4I6X9 U13357 ( .A(n688), .B(n686), .C(n673), .D(n5171), .Z(n5564)
         );
  HS65_LL_AOI222X2 U13358 ( .A(n689), .B(n670), .C(n674), .D(n5582), .E(n684), 
        .F(n678), .Z(n5566) );
  HS65_LL_CBI4I1X5 U13359 ( .A(n4535), .B(n5579), .C(n5581), .D(n5583), .Z(
        n5565) );
  HS65_LL_NAND4ABX3 U13360 ( .A(n4020), .B(n4021), .C(n4022), .D(n4023), .Z(
        n2713) );
  HS65_LL_CB4I6X9 U13361 ( .A(n441), .B(n440), .C(n407), .D(n3861), .Z(n4020)
         );
  HS65_LL_CBI4I1X5 U13362 ( .A(n2998), .B(n3203), .C(n3396), .D(n4043), .Z(
        n4021) );
  HS65_LL_AOI222X2 U13363 ( .A(n418), .B(n439), .C(n405), .D(n4042), .E(n411), 
        .F(n443), .Z(n4022) );
  HS65_LL_NAND4ABX3 U13364 ( .A(n7131), .B(n7132), .C(n7133), .D(n7134), .Z(
        n2808) );
  HS65_LL_CBI4I1X5 U13365 ( .A(n6388), .B(n6088), .C(n6568), .D(n6992), .Z(
        n7131) );
  HS65_LL_AOI212X4 U13366 ( .A(n279), .B(n303), .C(n278), .D(n6099), .E(n7150), 
        .Z(n7133) );
  HS65_LL_CBI4I1X5 U13367 ( .A(n7151), .B(n6085), .C(n6196), .D(n7152), .Z(
        n7132) );
  HS65_LL_NAND4ABX3 U13368 ( .A(n5539), .B(n5540), .C(n5541), .D(n5542), .Z(
        n2816) );
  HS65_LL_CBI4I1X5 U13369 ( .A(n4795), .B(n4495), .C(n4975), .D(n5400), .Z(
        n5539) );
  HS65_LL_AOI212X4 U13370 ( .A(n454), .B(n478), .C(n453), .D(n4506), .E(n5558), 
        .Z(n5541) );
  HS65_LL_CBI4I1X5 U13371 ( .A(n5559), .B(n4492), .C(n4603), .D(n5560), .Z(
        n5540) );
  HS65_LL_NAND4ABX3 U13372 ( .A(n3914), .B(n3915), .C(n3916), .D(n3917), .Z(
        n2673) );
  HS65_LL_CB4I6X9 U13373 ( .A(n221), .B(n220), .C(n200), .D(n3507), .Z(n3914)
         );
  HS65_LL_CBI4I1X5 U13374 ( .A(n2861), .B(n2938), .C(n3114), .D(n3930), .Z(
        n3915) );
  HS65_LL_AOI222X2 U13375 ( .A(n193), .B(n213), .C(n201), .D(n3929), .E(n197), 
        .F(n218), .Z(n3916) );
  HS65_LL_NAND4ABX3 U13376 ( .A(n5611), .B(n5612), .C(n5613), .D(n5614), .Z(
        n2815) );
  HS65_LL_CB4I6X9 U13377 ( .A(n474), .B(n473), .C(n454), .D(n5402), .Z(n5611)
         );
  HS65_LL_AOI222X2 U13378 ( .A(n480), .B(n461), .C(n453), .D(n5636), .E(n475), 
        .F(n450), .Z(n5613) );
  HS65_LL_CBI4I1X5 U13379 ( .A(n4604), .B(n5554), .C(n5630), .D(n5637), .Z(
        n5612) );
  HS65_LL_NAND4ABX3 U13380 ( .A(n9053), .B(n9054), .C(n9055), .D(n9056), .Z(
        n2800) );
  HS65_LL_CBI4I1X5 U13381 ( .A(n7662), .B(n7870), .C(n8449), .D(n8790), .Z(
        n9053) );
  HS65_LL_AOI212X4 U13382 ( .A(n111), .B(n125), .C(n112), .D(n7880), .E(n9108), 
        .Z(n9055) );
  HS65_LL_CBI4I1X5 U13383 ( .A(n8809), .B(n7714), .C(n7724), .D(n9110), .Z(
        n9054) );
  HS65_LL_NOR4ABX2 U13384 ( .A(n8642), .B(n8483), .C(n8637), .D(n8938), .Z(
        n8937) );
  HS65_LL_OAI212X5 U13385 ( .A(n7971), .B(n7861), .C(n8238), .D(n8302), .E(
        n7754), .Z(n8938) );
  HS65_LL_NAND4ABX3 U13386 ( .A(n3953), .B(n3954), .C(n3955), .D(n3956), .Z(
        n2708) );
  HS65_LL_AOI212X4 U13387 ( .A(n437), .B(n407), .C(n405), .D(n2843), .E(n3971), 
        .Z(n3955) );
  HS65_LL_CBI4I1X5 U13388 ( .A(n3198), .B(n2831), .C(n2994), .D(n3868), .Z(
        n3953) );
  HS65_LL_CBI4I1X5 U13389 ( .A(n3973), .B(n2829), .C(n2997), .D(n3974), .Z(
        n3954) );
  HS65_LL_NAND2X7 U13390 ( .A(n4329), .B(n4330), .Z(n2830) );
  HS65_LL_NAND4ABX3 U13391 ( .A(n5668), .B(n5669), .C(n5670), .D(n5671), .Z(
        n3209) );
  HS65_LL_NOR4ABX2 U13392 ( .A(n5160), .B(n5672), .C(n5142), .D(n4631), .Z(
        n5671) );
  HS65_LL_MX41X7 U13393 ( .D0(n690), .S0(n4521), .D1(n665), .S1(n686), .D2(
        n669), .S2(n701), .D3(n688), .S3(n674), .Z(n5668) );
  HS65_LL_MX41X7 U13394 ( .D0(n692), .S0(n671), .D1(n702), .S1(n677), .D2(n678), .S2(n691), .D3(n672), .S3(n4638), .Z(n5669) );
  HS65_LL_NAND4ABX3 U13395 ( .A(n7260), .B(n7261), .C(n7262), .D(n7263), .Z(
        n3006) );
  HS65_LL_NOR4ABX2 U13396 ( .A(n6752), .B(n7264), .C(n6734), .D(n6224), .Z(
        n7263) );
  HS65_LL_MX41X7 U13397 ( .D0(n514), .S0(n6114), .D1(n489), .S1(n510), .D2(
        n493), .S2(n525), .D3(n512), .S3(n498), .Z(n7260) );
  HS65_LL_MX41X7 U13398 ( .D0(n516), .S0(n495), .D1(n526), .S1(n501), .D2(n502), .S2(n515), .D3(n496), .S3(n6231), .Z(n7261) );
  HS65_LL_NOR4ABX2 U13399 ( .A(n4488), .B(n4489), .C(n4490), .D(n4491), .Z(
        n2821) );
  HS65_LL_OAI212X5 U13400 ( .A(n4492), .B(n4493), .C(n4494), .D(n4495), .E(
        n4496), .Z(n4491) );
  HS65_LL_NAND4ABX3 U13401 ( .A(n4502), .B(n4503), .C(n4504), .D(n4505), .Z(
        n4490) );
  HS65_LL_AOI212X4 U13402 ( .A(n451), .B(n479), .C(n455), .D(n472), .E(n4507), 
        .Z(n4489) );
  HS65_LL_NOR4ABX2 U13403 ( .A(n6081), .B(n6082), .C(n6083), .D(n6084), .Z(
        n2813) );
  HS65_LL_OAI212X5 U13404 ( .A(n6085), .B(n6086), .C(n6087), .D(n6088), .E(
        n6089), .Z(n6084) );
  HS65_LL_NAND4ABX3 U13405 ( .A(n6095), .B(n6096), .C(n6097), .D(n6098), .Z(
        n6083) );
  HS65_LL_AOI212X4 U13406 ( .A(n276), .B(n304), .C(n280), .D(n297), .E(n6100), 
        .Z(n6082) );
  HS65_LL_NAND4ABX3 U13407 ( .A(n2902), .B(n2903), .C(n2904), .D(n2905), .Z(
        n2631) );
  HS65_LL_CBI4I1X5 U13408 ( .A(n2913), .B(n2914), .C(n2915), .D(n2916), .Z(
        n2903) );
  HS65_LL_CBI4I1X5 U13409 ( .A(n2917), .B(n2918), .C(n2919), .D(n2920), .Z(
        n2902) );
  HS65_LL_AOI212X4 U13410 ( .A(n149), .B(n178), .C(n154), .D(n174), .E(n2911), 
        .Z(n2904) );
  HS65_LL_IVX9 U13411 ( .A(n4712), .Z(n39) );
  HS65_LL_IVX9 U13412 ( .A(n6305), .Z(n561) );
  HS65_LL_IVX9 U13413 ( .A(n1519), .Z(n819) );
  HS65_LL_IVX9 U13414 ( .A(n2271), .Z(n901) );
  HS65_LL_IVX9 U13415 ( .A(n1143), .Z(n860) );
  HS65_LL_IVX9 U13416 ( .A(n1895), .Z(n778) );
  HS65_LL_NAND2X7 U13417 ( .A(n2587), .B(n2596), .Z(n2238) );
  HS65_LL_NAND2X7 U13418 ( .A(n1835), .B(n1844), .Z(n1486) );
  HS65_LL_NAND2X7 U13419 ( .A(n2211), .B(n2220), .Z(n1862) );
  HS65_LL_NAND2X7 U13420 ( .A(n1459), .B(n1468), .Z(n1110) );
  HS65_LL_NAND4ABX3 U13421 ( .A(n8934), .B(n8935), .C(n8936), .D(n8937), .Z(
        n2751) );
  HS65_LL_CBI4I1X5 U13422 ( .A(n7858), .B(n8649), .C(n7966), .D(n8271), .Z(
        n8934) );
  HS65_LL_AOI222X2 U13423 ( .A(n369), .B(n398), .C(n373), .D(n8993), .E(n395), 
        .F(n375), .Z(n8936) );
  HS65_LL_CBI4I1X5 U13424 ( .A(n7852), .B(n7860), .C(n7750), .D(n8994), .Z(
        n8935) );
  HS65_LL_IVX9 U13425 ( .A(n4485), .Z(n9) );
  HS65_LL_IVX9 U13426 ( .A(n6078), .Z(n531) );
  HS65_LL_IVX9 U13427 ( .A(n8397), .Z(n585) );
  HS65_LL_IVX9 U13428 ( .A(n8449), .Z(n105) );
  HS65_LL_IVX9 U13429 ( .A(n7662), .Z(n134) );
  HS65_LL_IVX9 U13430 ( .A(n7622), .Z(n614) );
  HS65_LL_IVX9 U13431 ( .A(n5502), .Z(n14) );
  HS65_LL_IVX9 U13432 ( .A(n7094), .Z(n536) );
  HS65_LL_IVX9 U13433 ( .A(n8661), .Z(n395) );
  HS65_LL_NOR4ABX2 U13434 ( .A(n2825), .B(n2826), .C(n2827), .D(n2828), .Z(
        n2749) );
  HS65_LL_NAND4ABX3 U13435 ( .A(n2839), .B(n2840), .C(n2841), .D(n2842), .Z(
        n2827) );
  HS65_LL_OAI212X5 U13436 ( .A(n2829), .B(n2830), .C(n2831), .D(n2832), .E(
        n2833), .Z(n2828) );
  HS65_LL_AOI212X4 U13437 ( .A(n413), .B(n438), .C(n406), .D(n435), .E(n2844), 
        .Z(n2826) );
  HS65_LL_NAND4ABX3 U13438 ( .A(n5878), .B(n5879), .C(n5880), .D(n5881), .Z(
        n2814) );
  HS65_LL_NOR4ABX2 U13439 ( .A(n5392), .B(n5882), .C(n5374), .D(n4777), .Z(
        n5881) );
  HS65_LL_MX41X7 U13440 ( .D0(n477), .S0(n4606), .D1(n462), .S1(n473), .D2(
        n458), .S2(n467), .D3(n474), .S3(n453), .Z(n5878) );
  HS65_LL_MX41X7 U13441 ( .D0(n478), .S0(n459), .D1(n469), .S1(n449), .D2(n450), .S2(n479), .D3(n460), .S3(n4784), .Z(n5879) );
  HS65_LL_NAND4ABX3 U13442 ( .A(n7470), .B(n7471), .C(n7472), .D(n7473), .Z(
        n2806) );
  HS65_LL_NOR4ABX2 U13443 ( .A(n6984), .B(n7474), .C(n6966), .D(n6370), .Z(
        n7473) );
  HS65_LL_MX41X7 U13444 ( .D0(n302), .S0(n6199), .D1(n287), .S1(n298), .D2(
        n283), .S2(n292), .D3(n299), .S3(n278), .Z(n7470) );
  HS65_LL_MX41X7 U13445 ( .D0(n303), .S0(n284), .D1(n294), .S1(n274), .D2(n275), .S2(n304), .D3(n285), .S3(n6377), .Z(n7471) );
  HS65_LL_NAND4ABX3 U13446 ( .A(n7704), .B(n7705), .C(n7706), .D(n7707), .Z(
        n2798) );
  HS65_LL_MX41X7 U13447 ( .D0(n125), .S0(n96), .D1(n108), .S1(n122), .D2(n106), 
        .S2(n126), .D3(n100), .S3(n7738), .Z(n7705) );
  HS65_LL_MX41X7 U13448 ( .D0(n127), .S0(n7737), .D1(n104), .S1(n137), .D2(n99), .S2(n123), .D3(n134), .S3(n112), .Z(n7704) );
  HS65_LL_NOR4ABX2 U13449 ( .A(n7708), .B(n7709), .C(n7710), .D(n7711), .Z(
        n7707) );
  HS65_LL_IVX9 U13450 ( .A(n8018), .Z(n135) );
  HS65_LL_IVX9 U13451 ( .A(n2881), .Z(n658) );
  HS65_LL_IVX9 U13452 ( .A(n4608), .Z(n475) );
  HS65_LL_IVX9 U13453 ( .A(n4591), .Z(n258) );
  HS65_LL_IVX9 U13454 ( .A(n6184), .Z(n73) );
  HS65_LL_IVX9 U13455 ( .A(n6201), .Z(n300) );
  HS65_LL_IVX9 U13456 ( .A(n6117), .Z(n508) );
  HS65_LL_IVX9 U13457 ( .A(n4524), .Z(n684) );
  HS65_LL_IVX9 U13458 ( .A(n7821), .Z(n592) );
  HS65_LL_IVX9 U13459 ( .A(n7919), .Z(n112) );
  HS65_LL_IVX9 U13460 ( .A(n3097), .Z(n209) );
  HS65_LL_IVX9 U13461 ( .A(n2829), .Z(n427) );
  HS65_LL_IVX9 U13462 ( .A(n3253), .Z(n172) );
  HS65_LL_IVX9 U13463 ( .A(n3464), .Z(n201) );
  HS65_LL_IVX9 U13464 ( .A(n2992), .Z(n405) );
  HS65_LL_IVX9 U13465 ( .A(n2981), .Z(n624) );
  HS65_LL_IVX9 U13466 ( .A(n8871), .Z(n353) );
  HS65_LL_IVX9 U13467 ( .A(n2291), .Z(n885) );
  HS65_LL_IVX9 U13468 ( .A(n1163), .Z(n844) );
  HS65_LL_IVX9 U13469 ( .A(n1915), .Z(n762) );
  HS65_LL_IVX9 U13470 ( .A(n4484), .Z(n29) );
  HS65_LL_IVX9 U13471 ( .A(n6077), .Z(n551) );
  HS65_LL_IVX9 U13472 ( .A(n4572), .Z(n33) );
  HS65_LL_IVX9 U13473 ( .A(n6165), .Z(n555) );
  HS65_LL_OAI212X5 U13474 ( .A(n2005), .B(n1882), .C(n1908), .D(n1870), .E(
        n2006), .Z(n1995) );
  HS65_LL_NOR2X6 U13475 ( .A(n790), .B(n779), .Z(n2005) );
  HS65_LL_OAI21X3 U13476 ( .A(n792), .B(n786), .C(n766), .Z(n2006) );
  HS65_LL_OAI212X5 U13477 ( .A(n1253), .B(n1130), .C(n1156), .D(n1118), .E(
        n1254), .Z(n1243) );
  HS65_LL_NOR2X6 U13478 ( .A(n872), .B(n861), .Z(n1253) );
  HS65_LL_OAI21X3 U13479 ( .A(n874), .B(n868), .C(n848), .Z(n1254) );
  HS65_LL_IVX9 U13480 ( .A(n1539), .Z(n803) );
  HS65_LL_NAND4ABX3 U13481 ( .A(n5517), .B(n5518), .C(n5519), .D(n5520), .Z(
        n2792) );
  HS65_LL_CBI4I1X5 U13482 ( .A(n4734), .B(n4456), .C(n4922), .D(n5285), .Z(
        n5517) );
  HS65_LL_AOI212X4 U13483 ( .A(n237), .B(n261), .C(n236), .D(n4467), .E(n5536), 
        .Z(n5519) );
  HS65_LL_CBI4I1X5 U13484 ( .A(n5537), .B(n4453), .C(n4586), .D(n5538), .Z(
        n5518) );
  HS65_LL_NAND4ABX3 U13485 ( .A(n7109), .B(n7110), .C(n7111), .D(n7112), .Z(
        n2784) );
  HS65_LL_CBI4I1X5 U13486 ( .A(n6349), .B(n6049), .C(n6515), .D(n6877), .Z(
        n7109) );
  HS65_LL_AOI212X4 U13487 ( .A(n58), .B(n85), .C(n59), .D(n6060), .E(n7128), 
        .Z(n7111) );
  HS65_LL_CBI4I1X5 U13488 ( .A(n7129), .B(n6046), .C(n6179), .D(n7130), .Z(
        n7110) );
  HS65_LL_IVX9 U13489 ( .A(n1116), .Z(n868) );
  HS65_LL_IVX9 U13490 ( .A(n1868), .Z(n786) );
  HS65_LL_IVX9 U13491 ( .A(n3280), .Z(n178) );
  HS65_LL_IVX9 U13492 ( .A(n7940), .Z(n355) );
  HS65_LL_IVX9 U13493 ( .A(n3135), .Z(n650) );
  HS65_LL_IVX9 U13494 ( .A(n3048), .Z(n166) );
  HS65_LL_IVX9 U13495 ( .A(n8421), .Z(n616) );
  HS65_LL_IVX9 U13496 ( .A(n8473), .Z(n136) );
  HS65_LL_IVX9 U13497 ( .A(n5588), .Z(n241) );
  HS65_LL_IVX9 U13498 ( .A(n5630), .Z(n458) );
  HS65_LL_IVX9 U13499 ( .A(n7180), .Z(n57) );
  HS65_LL_IVX9 U13500 ( .A(n7222), .Z(n283) );
  HS65_LL_IVX9 U13501 ( .A(n7173), .Z(n493) );
  HS65_LL_IVX9 U13502 ( .A(n5581), .Z(n669) );
  HS65_LL_IVX9 U13503 ( .A(n1492), .Z(n827) );
  HS65_LL_IVX9 U13504 ( .A(n2244), .Z(n909) );
  HS65_LL_IVX9 U13505 ( .A(n7751), .Z(n390) );
  HS65_LL_IVX9 U13506 ( .A(n4734), .Z(n257) );
  HS65_LL_IVX9 U13507 ( .A(n4795), .Z(n474) );
  HS65_LL_IVX9 U13508 ( .A(n6349), .Z(n76) );
  HS65_LL_IVX9 U13509 ( .A(n6388), .Z(n299) );
  HS65_LL_IVX9 U13510 ( .A(n6242), .Z(n512) );
  HS65_LL_IVX9 U13511 ( .A(n4649), .Z(n688) );
  HS65_LL_IVX9 U13512 ( .A(n3588), .Z(n156) );
  HS65_LL_IVX9 U13513 ( .A(n3475), .Z(n188) );
  HS65_LL_IVX9 U13514 ( .A(n3972), .Z(n443) );
  HS65_LL_IVX9 U13515 ( .A(n6254), .Z(n567) );
  HS65_LL_IVX9 U13516 ( .A(n4661), .Z(n45) );
  HS65_LL_NAND2X7 U13517 ( .A(n8925), .B(n8918), .Z(n7952) );
  HS65_LL_NOR4ABX2 U13518 ( .A(n4577), .B(n4578), .C(n4579), .D(n4580), .Z(
        n2796) );
  HS65_LL_CBI4I6X5 U13519 ( .A(n234), .B(n4589), .C(n259), .D(n4590), .Z(n4578) );
  HS65_LL_CBI4I1X5 U13520 ( .A(n4586), .B(n4454), .C(n4587), .D(n4588), .Z(
        n4579) );
  HS65_LL_AOI212X4 U13521 ( .A(n253), .B(n243), .C(n267), .D(n235), .E(n4592), 
        .Z(n4577) );
  HS65_LL_NOR4ABX2 U13522 ( .A(n6170), .B(n6171), .C(n6172), .D(n6173), .Z(
        n2788) );
  HS65_LL_CBI4I6X5 U13523 ( .A(n63), .B(n6182), .C(n77), .D(n6183), .Z(n6171)
         );
  HS65_LL_CBI4I1X5 U13524 ( .A(n6179), .B(n6047), .C(n6180), .D(n6181), .Z(
        n6172) );
  HS65_LL_AOI212X4 U13525 ( .A(n88), .B(n56), .C(n81), .D(n66), .E(n6185), .Z(
        n6170) );
  HS65_LL_IVX9 U13526 ( .A(n3198), .Z(n441) );
  HS65_LL_IVX9 U13527 ( .A(n4453), .Z(n268) );
  HS65_LL_IVX9 U13528 ( .A(n4492), .Z(n485) );
  HS65_LL_IVX9 U13529 ( .A(n6046), .Z(n82) );
  HS65_LL_IVX9 U13530 ( .A(n6085), .Z(n310) );
  HS65_LL_IVX9 U13531 ( .A(n6443), .Z(n518) );
  HS65_LL_IVX9 U13532 ( .A(n4850), .Z(n694) );
  HS65_LL_IVX9 U13533 ( .A(n3952), .Z(n652) );
  HS65_LL_NAND4ABX3 U13534 ( .A(n4442), .B(n4443), .C(n4444), .D(n4445), .Z(
        n2797) );
  HS65_LL_OAI212X5 U13535 ( .A(n4453), .B(n4454), .C(n4455), .D(n4456), .E(
        n4457), .Z(n4443) );
  HS65_LL_NAND4ABX3 U13536 ( .A(n4463), .B(n4464), .C(n4465), .D(n4466), .Z(
        n4442) );
  HS65_LL_AOI212X4 U13537 ( .A(n234), .B(n262), .C(n238), .D(n255), .E(n4446), 
        .Z(n4445) );
  HS65_LL_NAND4ABX3 U13538 ( .A(n6035), .B(n6036), .C(n6037), .D(n6038), .Z(
        n2789) );
  HS65_LL_OAI212X5 U13539 ( .A(n6046), .B(n6047), .C(n6048), .D(n6049), .E(
        n6050), .Z(n6036) );
  HS65_LL_NAND4ABX3 U13540 ( .A(n6056), .B(n6057), .C(n6058), .D(n6059), .Z(
        n6035) );
  HS65_LL_AOI212X4 U13541 ( .A(n63), .B(n84), .C(n60), .D(n90), .E(n6039), .Z(
        n6038) );
  HS65_LL_NAND4ABX3 U13542 ( .A(n3350), .B(n3351), .C(n3352), .D(n3353), .Z(
        n2698) );
  HS65_LL_NAND4ABX3 U13543 ( .A(n3408), .B(n3409), .C(n3410), .D(n3411), .Z(
        n3350) );
  HS65_LL_OAI212X5 U13544 ( .A(n3404), .B(n2832), .C(n3405), .D(n3406), .E(
        n3407), .Z(n3351) );
  HS65_LL_AOI212X4 U13545 ( .A(n405), .B(n426), .C(n432), .D(n409), .E(n3354), 
        .Z(n3353) );
  HS65_LL_IVX9 U13546 ( .A(n3928), .Z(n218) );
  HS65_LL_IVX9 U13547 ( .A(n4668), .Z(n30) );
  HS65_LL_IVX9 U13548 ( .A(n6261), .Z(n552) );
  HS65_LL_IVX9 U13549 ( .A(n5013), .Z(n19) );
  HS65_LL_IVX9 U13550 ( .A(n6606), .Z(n541) );
  HS65_LL_IVX9 U13551 ( .A(n2933), .Z(n221) );
  HS65_LL_IVX9 U13552 ( .A(n7858), .Z(n393) );
  HS65_LL_IVX9 U13553 ( .A(n7636), .Z(n600) );
  HS65_LL_IVX9 U13554 ( .A(n7657), .Z(n120) );
  HS65_LL_IVX9 U13555 ( .A(n6455), .Z(n524) );
  HS65_LL_IVX9 U13556 ( .A(n4862), .Z(n700) );
  HS65_LL_IVX9 U13557 ( .A(n4876), .Z(n253) );
  HS65_LL_IVX9 U13558 ( .A(n6581), .Z(n295) );
  HS65_LL_IVX9 U13559 ( .A(n6469), .Z(n88) );
  HS65_LL_IVX9 U13560 ( .A(n4988), .Z(n470) );
  HS65_LL_IVX9 U13561 ( .A(n3293), .Z(n646) );
  HS65_LL_NAND4ABX3 U13562 ( .A(n6526), .B(n6527), .C(n6528), .D(n6529), .Z(
        n2810) );
  HS65_LL_NAND4ABX3 U13563 ( .A(n6583), .B(n6584), .C(n6585), .D(n6586), .Z(
        n6526) );
  HS65_LL_OAI212X5 U13564 ( .A(n6579), .B(n6087), .C(n6580), .D(n6581), .E(
        n6582), .Z(n6527) );
  HS65_LL_AOI212X4 U13565 ( .A(n278), .B(n308), .C(n294), .D(n274), .E(n6530), 
        .Z(n6529) );
  HS65_LL_NAND4ABX3 U13566 ( .A(n4933), .B(n4934), .C(n4935), .D(n4936), .Z(
        n2818) );
  HS65_LL_NAND4ABX3 U13567 ( .A(n4990), .B(n4991), .C(n4992), .D(n4993), .Z(
        n4933) );
  HS65_LL_OAI212X5 U13568 ( .A(n4986), .B(n4494), .C(n4987), .D(n4988), .E(
        n4989), .Z(n4934) );
  HS65_LL_AOI212X4 U13569 ( .A(n453), .B(n483), .C(n469), .D(n449), .E(n4937), 
        .Z(n4936) );
  HS65_LL_IVX9 U13570 ( .A(n2146), .Z(n758) );
  HS65_LL_IVX9 U13571 ( .A(n1745), .Z(n824) );
  HS65_LL_IVX9 U13572 ( .A(n8357), .Z(n340) );
  HS65_LL_IVX9 U13573 ( .A(n1394), .Z(n840) );
  HS65_LL_IVX9 U13574 ( .A(n1770), .Z(n799) );
  HS65_LL_IVX9 U13575 ( .A(n2522), .Z(n881) );
  HS65_LL_IVX9 U13576 ( .A(n2497), .Z(n906) );
  HS65_LL_IVX9 U13577 ( .A(n1369), .Z(n865) );
  HS65_LL_IVX9 U13578 ( .A(n2121), .Z(n783) );
  HS65_LL_IVX9 U13579 ( .A(n7783), .Z(n610) );
  HS65_LL_IVX9 U13580 ( .A(n7882), .Z(n130) );
  HS65_LL_NAND4ABX3 U13581 ( .A(n7932), .B(n7933), .C(n7934), .D(n7935), .Z(
        n3004) );
  HS65_LL_CBI4I1X5 U13582 ( .A(n7951), .B(n7952), .C(n7953), .D(n321), .Z(
        n7932) );
  HS65_LL_CBI4I1X5 U13583 ( .A(n7947), .B(n7948), .C(n7949), .D(n7950), .Z(
        n7933) );
  HS65_LL_AOI212X4 U13584 ( .A(n345), .B(n334), .C(n328), .D(n340), .E(n7945), 
        .Z(n7934) );
  HS65_LL_OAI212X5 U13585 ( .A(n7918), .B(n7652), .C(n7919), .D(n7920), .E(
        n7921), .Z(n7917) );
  HS65_LL_NOR3X4 U13586 ( .A(n119), .B(n124), .C(n123), .Z(n7918) );
  HS65_LL_OAI21X3 U13587 ( .A(n105), .B(n100), .C(n131), .Z(n7921) );
  HS65_LL_IVX9 U13588 ( .A(n3994), .Z(n169) );
  HS65_LL_NOR4ABX2 U13589 ( .A(n5584), .B(n5585), .C(n5586), .D(n5587), .Z(
        n2791) );
  HS65_LL_CB4I6X9 U13590 ( .A(n257), .B(n256), .C(n237), .D(n5287), .Z(n5586)
         );
  HS65_LL_AOI222X2 U13591 ( .A(n263), .B(n244), .C(n236), .D(n5610), .E(n258), 
        .F(n233), .Z(n5584) );
  HS65_LL_CBI4I1X5 U13592 ( .A(n4587), .B(n5532), .C(n5588), .D(n5589), .Z(
        n5587) );
  HS65_LL_NOR4ABX2 U13593 ( .A(n7176), .B(n7177), .C(n7178), .D(n7179), .Z(
        n2783) );
  HS65_LL_CB4I6X9 U13594 ( .A(n76), .B(n74), .C(n58), .D(n6879), .Z(n7178) );
  HS65_LL_AOI222X2 U13595 ( .A(n86), .B(n55), .C(n59), .D(n7202), .E(n73), .F(
        n64), .Z(n7176) );
  HS65_LL_CBI4I1X5 U13596 ( .A(n6180), .B(n7124), .C(n7180), .D(n7181), .Z(
        n7179) );
  HS65_LL_NOR4ABX2 U13597 ( .A(n7614), .B(n7615), .C(n7616), .D(n7617), .Z(
        n2775) );
  HS65_LL_CBI4I1X5 U13598 ( .A(n7622), .B(n7623), .C(n7624), .D(n7625), .Z(
        n7616) );
  HS65_LL_CBI4I1X5 U13599 ( .A(n7618), .B(n7619), .C(n7620), .D(n7621), .Z(
        n7617) );
  HS65_LL_AOI222X2 U13600 ( .A(n604), .B(n578), .C(n592), .D(n7635), .E(n615), 
        .F(n586), .Z(n7614) );
  HS65_LL_IVX9 U13601 ( .A(n8082), .Z(n389) );
  HS65_LL_IVX9 U13602 ( .A(n1524), .Z(n826) );
  HS65_LL_IVX9 U13603 ( .A(n2276), .Z(n908) );
  HS65_LL_IVX9 U13604 ( .A(n1148), .Z(n867) );
  HS65_LL_IVX9 U13605 ( .A(n1900), .Z(n785) );
  HS65_LL_IVX9 U13606 ( .A(n6278), .Z(n563) );
  HS65_LL_IVX9 U13607 ( .A(n4685), .Z(n41) );
  HS65_LL_OAI212X5 U13608 ( .A(n8965), .B(n8238), .C(n7993), .D(n8207), .E(
        n8966), .Z(n8964) );
  HS65_LL_OAI21X3 U13609 ( .A(n378), .B(n370), .C(n391), .Z(n8966) );
  HS65_LL_NOR3X4 U13610 ( .A(n398), .B(n386), .C(n387), .Z(n8965) );
  HS65_LL_NAND4ABX3 U13611 ( .A(n6110), .B(n6111), .C(n6112), .D(n6113), .Z(
        n3207) );
  HS65_LL_CBI4I6X5 U13612 ( .A(n503), .B(n6114), .C(n509), .D(n6115), .Z(n6113) );
  HS65_LL_CBI4I1X5 U13613 ( .A(n6126), .B(n6127), .C(n6128), .D(n6129), .Z(
        n6110) );
  HS65_LL_AOI212X4 U13614 ( .A(n524), .B(n496), .C(n520), .D(n504), .E(n6119), 
        .Z(n6112) );
  HS65_LL_NAND4ABX3 U13615 ( .A(n4517), .B(n4518), .C(n4519), .D(n4520), .Z(
        n3532) );
  HS65_LL_CBI4I6X5 U13616 ( .A(n679), .B(n4521), .C(n685), .D(n4522), .Z(n4520) );
  HS65_LL_CBI4I1X5 U13617 ( .A(n4533), .B(n4534), .C(n4535), .D(n4536), .Z(
        n4517) );
  HS65_LL_AOI212X4 U13618 ( .A(n700), .B(n672), .C(n696), .D(n680), .E(n4526), 
        .Z(n4519) );
  HS65_LL_IVX9 U13619 ( .A(n8339), .Z(n349) );
  HS65_LL_NAND2X7 U13620 ( .A(n3133), .B(n2889), .Z(n3311) );
  HS65_LL_IVX9 U13621 ( .A(n7631), .Z(n607) );
  HS65_LL_IVX9 U13622 ( .A(n7651), .Z(n127) );
  HS65_LL_IVX9 U13623 ( .A(n3112), .Z(n212) );
  HS65_LL_IVX9 U13624 ( .A(n4549), .Z(n37) );
  HS65_LL_IVX9 U13625 ( .A(n6142), .Z(n559) );
  HS65_LL_IVX9 U13626 ( .A(n2520), .Z(n890) );
  HS65_LL_IVX9 U13627 ( .A(n8067), .Z(n391) );
  HS65_LL_IVX9 U13628 ( .A(n4593), .Z(n236) );
  HS65_LL_IVX9 U13629 ( .A(n4610), .Z(n453) );
  HS65_LL_IVX9 U13630 ( .A(n6186), .Z(n59) );
  HS65_LL_IVX9 U13631 ( .A(n6203), .Z(n278) );
  HS65_LL_IVX9 U13632 ( .A(n2144), .Z(n767) );
  HS65_LL_IVX9 U13633 ( .A(n1392), .Z(n849) );
  HS65_LL_IVX9 U13634 ( .A(n1768), .Z(n808) );
  HS65_LL_NOR2X6 U13635 ( .A(n3950), .B(n3133), .Z(n3742) );
  HS65_LL_IVX9 U13636 ( .A(n7951), .Z(n325) );
  HS65_LL_IVX9 U13637 ( .A(n7993), .Z(n397) );
  HS65_LL_IVX9 U13638 ( .A(n5265), .Z(n262) );
  HS65_LL_IVX9 U13639 ( .A(n5380), .Z(n479) );
  HS65_LL_IVX9 U13640 ( .A(n6972), .Z(n304) );
  HS65_LL_IVX9 U13641 ( .A(n6740), .Z(n515) );
  HS65_LL_IVX9 U13642 ( .A(n6857), .Z(n84) );
  HS65_LL_IVX9 U13643 ( .A(n2876), .Z(n659) );
  HS65_LL_IVX9 U13644 ( .A(n3926), .Z(n220) );
  HS65_LL_IVX9 U13645 ( .A(n3970), .Z(n440) );
  HS65_LL_IVX9 U13646 ( .A(n7653), .Z(n132) );
  HS65_LL_IVX9 U13647 ( .A(n7633), .Z(n612) );
  HS65_LL_NAND2X7 U13648 ( .A(n9043), .B(n9020), .Z(n7806) );
  HS65_LL_NAND2X7 U13649 ( .A(n9101), .B(n9078), .Z(n7869) );
  HS65_LL_NOR2X6 U13650 ( .A(n8649), .B(n7965), .Z(n8264) );
  HS65_LL_IVX9 U13651 ( .A(n4500), .Z(n461) );
  HS65_LL_IVX9 U13652 ( .A(n6093), .Z(n286) );
  HS65_LL_IVX9 U13653 ( .A(n4461), .Z(n244) );
  HS65_LL_IVX9 U13654 ( .A(n6054), .Z(n55) );
  HS65_LL_IVX9 U13655 ( .A(n7088), .Z(n494) );
  HS65_LL_IVX9 U13656 ( .A(n5496), .Z(n670) );
  HS65_LL_IVX9 U13657 ( .A(n7850), .Z(n374) );
  HS65_LL_IVX9 U13658 ( .A(n2069), .Z(n763) );
  HS65_LL_IVX9 U13659 ( .A(n1317), .Z(n845) );
  HS65_LL_IVX9 U13660 ( .A(n3450), .Z(n211) );
  HS65_LL_IVX9 U13661 ( .A(n3035), .Z(n155) );
  HS65_LL_IVX9 U13662 ( .A(n2297), .Z(n889) );
  HS65_LL_IVX9 U13663 ( .A(n3950), .Z(n649) );
  HS65_LL_IVX9 U13664 ( .A(n8313), .Z(n341) );
  HS65_LL_IVX9 U13665 ( .A(n1162), .Z(n871) );
  HS65_LL_IVX9 U13666 ( .A(n1914), .Z(n789) );
  HS65_LL_IVX9 U13667 ( .A(n2445), .Z(n886) );
  HS65_LL_IVX9 U13668 ( .A(n6247), .Z(n520) );
  HS65_LL_IVX9 U13669 ( .A(n4654), .Z(n696) );
  HS65_LL_IVX9 U13670 ( .A(n4447), .Z(n267) );
  HS65_LL_IVX9 U13671 ( .A(n6101), .Z(n309) );
  HS65_LL_IVX9 U13672 ( .A(n6040), .Z(n81) );
  HS65_LL_IVX9 U13673 ( .A(n4508), .Z(n484) );
  HS65_LL_IVX9 U13674 ( .A(n8527), .Z(n343) );
  HS65_LL_IVX9 U13675 ( .A(n1921), .Z(n766) );
  HS65_LL_IVX9 U13676 ( .A(n1169), .Z(n848) );
  HS65_LL_IVX9 U13677 ( .A(n3184), .Z(n407) );
  HS65_LL_IVX9 U13678 ( .A(n1693), .Z(n804) );
  HS65_LL_IVX9 U13679 ( .A(n7183), .Z(n78) );
  HS65_LL_IVX9 U13680 ( .A(n5591), .Z(n264) );
  HS65_LL_IVX9 U13681 ( .A(n5616), .Z(n481) );
  HS65_LL_IVX9 U13682 ( .A(n7208), .Z(n306) );
  HS65_LL_IVX9 U13683 ( .A(n7164), .Z(n521) );
  HS65_LL_IVX9 U13684 ( .A(n1545), .Z(n807) );
  HS65_LL_IVX9 U13685 ( .A(n8302), .Z(n392) );
  HS65_LL_IVX9 U13686 ( .A(n1538), .Z(n830) );
  HS65_LL_IVX9 U13687 ( .A(n2290), .Z(n912) );
  HS65_LL_NOR2X6 U13688 ( .A(n2883), .B(n3133), .Z(n3672) );
  HS65_LL_IVX9 U13689 ( .A(n5508), .Z(n42) );
  HS65_LL_IVX9 U13690 ( .A(n7100), .Z(n564) );
  HS65_LL_IVX9 U13691 ( .A(n3397), .Z(n438) );
  HS65_LL_NOR2X6 U13692 ( .A(n7147), .B(n7222), .Z(n7052) );
  HS65_LL_NOR2X6 U13693 ( .A(n5533), .B(n5588), .Z(n5345) );
  HS65_LL_NOR2X6 U13694 ( .A(n7125), .B(n7180), .Z(n6937) );
  HS65_LL_IVX9 U13695 ( .A(n3343), .Z(n655) );
  HS65_LL_IVX9 U13696 ( .A(n2932), .Z(n200) );
  HS65_LL_IVX9 U13697 ( .A(n2838), .Z(n429) );
  HS65_LL_IVX9 U13698 ( .A(n3069), .Z(n210) );
  HS65_LL_IVX9 U13699 ( .A(n2846), .Z(n428) );
  HS65_LL_IVX9 U13700 ( .A(n2939), .Z(n216) );
  HS65_LL_NOR2X6 U13701 ( .A(n8178), .B(n7657), .Z(n8436) );
  HS65_LL_NOR2X6 U13702 ( .A(n7846), .B(n8082), .Z(n8075) );
  HS65_LL_IVX9 U13703 ( .A(n3134), .Z(n626) );
  HS65_LL_IVX9 U13704 ( .A(n5604), .Z(n256) );
  HS65_LL_IVX9 U13705 ( .A(n5629), .Z(n473) );
  HS65_LL_IVX9 U13706 ( .A(n7196), .Z(n74) );
  HS65_LL_IVX9 U13707 ( .A(n7221), .Z(n298) );
  HS65_LL_NOR2X6 U13708 ( .A(n2239), .B(n2276), .Z(n2461) );
  HS65_LL_NOR2X6 U13709 ( .A(n1487), .B(n1524), .Z(n1709) );
  HS65_LL_NOR2X6 U13710 ( .A(n1863), .B(n1900), .Z(n2085) );
  HS65_LL_NOR2X6 U13711 ( .A(n1111), .B(n1148), .Z(n1333) );
  HS65_LL_IVX9 U13712 ( .A(n3115), .Z(n214) );
  HS65_LL_NOR2X6 U13713 ( .A(n2970), .B(n3133), .Z(n3770) );
  HS65_LL_IVX9 U13714 ( .A(n4775), .Z(n454) );
  HS65_LL_IVX9 U13715 ( .A(n4733), .Z(n237) );
  HS65_LL_IVX9 U13716 ( .A(n6368), .Z(n279) );
  HS65_LL_IVX9 U13717 ( .A(n6329), .Z(n58) );
  HS65_LL_IVX9 U13718 ( .A(n6222), .Z(n497) );
  HS65_LL_IVX9 U13719 ( .A(n4629), .Z(n673) );
  HS65_LL_NOR2X6 U13720 ( .A(n7870), .B(n8183), .Z(n8820) );
  HS65_LL_NOR2X6 U13721 ( .A(n7831), .B(n8132), .Z(n8730) );
  HS65_LL_IVX9 U13722 ( .A(n7966), .Z(n371) );
  HS65_LL_IVX9 U13723 ( .A(n2258), .Z(n892) );
  HS65_LL_IVX9 U13724 ( .A(n2890), .Z(n660) );
  HS65_LL_IVX9 U13725 ( .A(n1882), .Z(n769) );
  HS65_LL_IVX9 U13726 ( .A(n1130), .Z(n851) );
  HS65_LL_IVX9 U13727 ( .A(n1532), .Z(n832) );
  HS65_LL_IVX9 U13728 ( .A(n3192), .Z(n417) );
  HS65_LL_IVX9 U13729 ( .A(n2926), .Z(n194) );
  HS65_LL_NOR2X6 U13730 ( .A(n2890), .B(n2981), .Z(n3744) );
  HS65_LL_IVX9 U13731 ( .A(n1506), .Z(n810) );
  HS65_LL_IVX9 U13732 ( .A(n4550), .Z(n10) );
  HS65_LL_IVX9 U13733 ( .A(n6143), .Z(n532) );
  HS65_LL_IVX9 U13734 ( .A(n2284), .Z(n914) );
  HS65_LL_IVX9 U13735 ( .A(n1156), .Z(n873) );
  HS65_LL_IVX9 U13736 ( .A(n1908), .Z(n791) );
  HS65_LL_IVX9 U13737 ( .A(n3224), .Z(n173) );
  HS65_LL_NOR2X6 U13738 ( .A(n4727), .B(n5591), .Z(n4916) );
  HS65_LL_NOR2X6 U13739 ( .A(n4789), .B(n5616), .Z(n4969) );
  HS65_LL_NOR2X6 U13740 ( .A(n6382), .B(n7208), .Z(n6562) );
  HS65_LL_NOR2X6 U13741 ( .A(n6343), .B(n7183), .Z(n6509) );
  HS65_LL_IVX9 U13742 ( .A(n8034), .Z(n324) );
  HS65_LL_IVX9 U13743 ( .A(n3054), .Z(n174) );
  HS65_LL_IVX9 U13744 ( .A(n4790), .Z(n472) );
  HS65_LL_IVX9 U13745 ( .A(n4728), .Z(n255) );
  HS65_LL_IVX9 U13746 ( .A(n6383), .Z(n297) );
  HS65_LL_IVX9 U13747 ( .A(n4644), .Z(n699) );
  HS65_LL_IVX9 U13748 ( .A(n6237), .Z(n523) );
  HS65_LL_IVX9 U13749 ( .A(n6344), .Z(n90) );
  HS65_LL_IVX9 U13750 ( .A(n4455), .Z(n247) );
  HS65_LL_IVX9 U13751 ( .A(n4494), .Z(n464) );
  HS65_LL_IVX9 U13752 ( .A(n6048), .Z(n68) );
  HS65_LL_IVX9 U13753 ( .A(n6087), .Z(n289) );
  HS65_LL_IVX9 U13754 ( .A(n6219), .Z(n490) );
  HS65_LL_IVX9 U13755 ( .A(n4626), .Z(n666) );
  HS65_LL_IVX9 U13756 ( .A(n4552), .Z(n18) );
  HS65_LL_IVX9 U13757 ( .A(n6145), .Z(n540) );
  HS65_LL_IVX9 U13758 ( .A(n8128), .Z(n580) );
  HS65_LL_IVX9 U13759 ( .A(n8179), .Z(n100) );
  HS65_LL_IVX9 U13760 ( .A(n7875), .Z(n131) );
  HS65_LL_IVX9 U13761 ( .A(n7836), .Z(n611) );
  HS65_LL_IVX9 U13762 ( .A(n3128), .Z(n635) );
  HS65_LL_IVX9 U13763 ( .A(n8028), .Z(n334) );
  HS65_LL_IVX9 U13764 ( .A(n5514), .Z(n31) );
  HS65_LL_IVX9 U13765 ( .A(n7106), .Z(n553) );
  HS65_LL_NOR2X6 U13766 ( .A(n4727), .B(n5265), .Z(n5342) );
  HS65_LL_NOR2X6 U13767 ( .A(n6382), .B(n6972), .Z(n7049) );
  HS65_LL_NOR2X6 U13768 ( .A(n6343), .B(n6857), .Z(n6934) );
  HS65_LL_IVX9 U13769 ( .A(n7960), .Z(n370) );
  HS65_LL_NOR2X6 U13770 ( .A(n7947), .B(n8357), .Z(n8360) );
  HS65_LL_IVX9 U13771 ( .A(n3204), .Z(n436) );
  HS65_LL_IVX9 U13772 ( .A(n6055), .Z(n79) );
  HS65_LL_IVX9 U13773 ( .A(n4462), .Z(n265) );
  HS65_LL_IVX9 U13774 ( .A(n4501), .Z(n482) );
  HS65_LL_IVX9 U13775 ( .A(n4523), .Z(n695) );
  HS65_LL_IVX9 U13776 ( .A(n4483), .Z(n40) );
  HS65_LL_IVX9 U13777 ( .A(n6094), .Z(n307) );
  HS65_LL_IVX9 U13778 ( .A(n6116), .Z(n519) );
  HS65_LL_IVX9 U13779 ( .A(n6076), .Z(n562) );
  HS65_LL_IVX9 U13780 ( .A(n2240), .Z(n916) );
  HS65_LL_IVX9 U13781 ( .A(n1488), .Z(n834) );
  HS65_LL_IVX9 U13782 ( .A(n1864), .Z(n793) );
  HS65_LL_IVX9 U13783 ( .A(n1112), .Z(n875) );
  HS65_LL_NOR2X6 U13784 ( .A(n1743), .B(n1532), .Z(n1607) );
  HS65_LL_NOR2X6 U13785 ( .A(n2246), .B(n2271), .Z(n2460) );
  HS65_LL_NOR2X6 U13786 ( .A(n1494), .B(n1519), .Z(n1708) );
  HS65_LL_NOR2X6 U13787 ( .A(n1870), .B(n1895), .Z(n2084) );
  HS65_LL_NOR2X6 U13788 ( .A(n1118), .B(n1143), .Z(n1332) );
  HS65_LL_IVX9 U13789 ( .A(n7650), .Z(n103) );
  HS65_LL_IVX9 U13790 ( .A(n7630), .Z(n583) );
  HS65_LL_IVX9 U13791 ( .A(n4732), .Z(n242) );
  HS65_LL_IVX9 U13792 ( .A(n4794), .Z(n459) );
  HS65_LL_IVX9 U13793 ( .A(n4648), .Z(n671) );
  HS65_LL_IVX9 U13794 ( .A(n6348), .Z(n54) );
  HS65_LL_IVX9 U13795 ( .A(n6387), .Z(n284) );
  HS65_LL_IVX9 U13796 ( .A(n6241), .Z(n495) );
  HS65_LL_IVX9 U13797 ( .A(n7961), .Z(n386) );
  HS65_LL_IVX9 U13798 ( .A(n8029), .Z(n347) );
  HS65_LL_NOR2X6 U13799 ( .A(n2495), .B(n2284), .Z(n2359) );
  HS65_LL_NOR2X6 U13800 ( .A(n2119), .B(n1908), .Z(n1983) );
  HS65_LL_NOR2X6 U13801 ( .A(n1367), .B(n1156), .Z(n1231) );
  HS65_LL_IVX9 U13802 ( .A(n2956), .Z(n189) );
  HS65_LL_NOR2X6 U13803 ( .A(n1487), .B(n1532), .Z(n1733) );
  HS65_LL_NOR2X6 U13804 ( .A(n8302), .B(n7960), .Z(n8105) );
  HS65_LL_NOR2X6 U13805 ( .A(n2831), .B(n3192), .Z(n3884) );
  HS65_LL_IVX9 U13806 ( .A(n4567), .Z(n44) );
  HS65_LL_IVX9 U13807 ( .A(n6160), .Z(n566) );
  HS65_LL_NOR2X6 U13808 ( .A(n2837), .B(n3193), .Z(n3839) );
  HS65_LL_NOR2X6 U13809 ( .A(n3116), .B(n2927), .Z(n3484) );
  HS65_LL_NOR2X6 U13810 ( .A(n2239), .B(n2284), .Z(n2485) );
  HS65_LL_NOR2X6 U13811 ( .A(n1111), .B(n1156), .Z(n1357) );
  HS65_LL_NOR2X6 U13812 ( .A(n1863), .B(n1908), .Z(n2109) );
  HS65_LL_IVX9 U13813 ( .A(n3042), .Z(n149) );
  HS65_LL_NOR2X6 U13814 ( .A(n1117), .B(n1157), .Z(n1311) );
  HS65_LL_NOR2X6 U13815 ( .A(n1869), .B(n1909), .Z(n2063) );
  HS65_LL_IVX9 U13816 ( .A(n4571), .Z(n16) );
  HS65_LL_IVX9 U13817 ( .A(n6164), .Z(n538) );
  HS65_LL_NOR2X6 U13818 ( .A(n2245), .B(n2285), .Z(n2439) );
  HS65_LL_NOR2X6 U13819 ( .A(n1493), .B(n1533), .Z(n1687) );
  HS65_LL_NOR2X6 U13820 ( .A(n2883), .B(n3128), .Z(n3769) );
  HS65_LL_IVX9 U13821 ( .A(n8057), .Z(n328) );
  HS65_LL_NOR2X6 U13822 ( .A(n2876), .B(n3134), .Z(n3762) );
  HS65_LL_IVX9 U13823 ( .A(n4643), .Z(n672) );
  HS65_LL_IVX9 U13824 ( .A(n6236), .Z(n496) );
  HS65_LL_IVX9 U13825 ( .A(n4727), .Z(n243) );
  HS65_LL_IVX9 U13826 ( .A(n6382), .Z(n285) );
  HS65_LL_IVX9 U13827 ( .A(n6343), .Z(n56) );
  HS65_LL_IVX9 U13828 ( .A(n4789), .Z(n460) );
  HS65_LL_NOR2X6 U13829 ( .A(n3203), .B(n3192), .Z(n3778) );
  HS65_LL_NOR2X6 U13830 ( .A(n8132), .B(n8421), .Z(n7690) );
  HS65_LL_NOR2X6 U13831 ( .A(n2889), .B(n3129), .Z(n3725) );
  HS65_LL_IVX9 U13832 ( .A(n2884), .Z(n640) );
  HS65_LL_IVX9 U13833 ( .A(n7965), .Z(n368) );
  HS65_LL_NOR2X6 U13834 ( .A(n7859), .B(n7961), .Z(n8247) );
  HS65_LL_IVX9 U13835 ( .A(n7905), .Z(n119) );
  HS65_LL_IVX9 U13836 ( .A(n7807), .Z(n599) );
  HS65_LL_IVX9 U13837 ( .A(n8033), .Z(n335) );
  HS65_LL_NOR2X6 U13838 ( .A(n1882), .B(n1914), .Z(n2102) );
  HS65_LL_NOR2X6 U13839 ( .A(n1130), .B(n1162), .Z(n1350) );
  HS65_LL_IVX9 U13840 ( .A(n1157), .Z(n850) );
  HS65_LL_IVX9 U13841 ( .A(n1909), .Z(n768) );
  HS65_LL_IVX9 U13842 ( .A(n2993), .Z(n419) );
  HS65_LL_IVX9 U13843 ( .A(n2968), .Z(n637) );
  HS65_LL_NOR2X6 U13844 ( .A(n2846), .B(n3184), .Z(n3877) );
  HS65_LL_IVX9 U13845 ( .A(n2285), .Z(n891) );
  HS65_LL_NOR2X6 U13846 ( .A(n2258), .B(n2290), .Z(n2478) );
  HS65_LL_NOR2X6 U13847 ( .A(n1506), .B(n1538), .Z(n1726) );
  HS65_LL_IVX9 U13848 ( .A(n1533), .Z(n809) );
  HS65_LL_NOR2X6 U13849 ( .A(n7750), .B(n8302), .Z(n8206) );
  HS65_LL_NOR2X6 U13850 ( .A(n2246), .B(n2333), .Z(n2482) );
  HS65_LL_NOR2X6 U13851 ( .A(n1118), .B(n1205), .Z(n1354) );
  HS65_LL_NOR2X6 U13852 ( .A(n1494), .B(n1581), .Z(n1730) );
  HS65_LL_NOR2X6 U13853 ( .A(n1870), .B(n1957), .Z(n2106) );
  HS65_LL_NOR2X6 U13854 ( .A(n2838), .B(n3412), .Z(n3881) );
  HS65_LL_NOR2X6 U13855 ( .A(n3069), .B(n3067), .Z(n3527) );
  HS65_LL_IVX9 U13856 ( .A(n1520), .Z(n823) );
  HS65_LL_IVX9 U13857 ( .A(n2272), .Z(n905) );
  HS65_LL_IVX9 U13858 ( .A(n1896), .Z(n782) );
  HS65_LL_IVX9 U13859 ( .A(n1144), .Z(n864) );
  HS65_LL_IVX9 U13860 ( .A(n8132), .Z(n576) );
  HS65_LL_IVX9 U13861 ( .A(n8183), .Z(n96) );
  HS65_LL_NOR2X6 U13862 ( .A(n8082), .B(n7847), .Z(n8222) );
  HS65_LL_IVX9 U13863 ( .A(n2855), .Z(n191) );
  HS65_LL_NOR2X6 U13864 ( .A(n2258), .B(n2273), .Z(n2399) );
  HS65_LL_IVX9 U13865 ( .A(n3193), .Z(n435) );
  HS65_LL_IVX9 U13866 ( .A(n2927), .Z(n223) );
  HS65_LL_NOR2X6 U13867 ( .A(n1882), .B(n1897), .Z(n2023) );
  HS65_LL_NOR2X6 U13868 ( .A(n1130), .B(n1145), .Z(n1271) );
  HS65_LL_IVX9 U13869 ( .A(n3133), .Z(n634) );
  HS65_LL_NOR2X6 U13870 ( .A(n1506), .B(n1521), .Z(n1647) );
  HS65_LL_NOR2X6 U13871 ( .A(n1914), .B(n1920), .Z(n2105) );
  HS65_LL_NOR2X6 U13872 ( .A(n1162), .B(n1168), .Z(n1353) );
  HS65_LL_NOR2X6 U13873 ( .A(n2846), .B(n2994), .Z(n3786) );
  HS65_LL_NOR2X6 U13874 ( .A(n3112), .B(n2856), .Z(n3428) );
  HS65_LL_NOR2X6 U13875 ( .A(n2290), .B(n2296), .Z(n2481) );
  HS65_LL_NOR2X6 U13876 ( .A(n8449), .B(n7882), .Z(n8815) );
  HS65_LL_NOR2X6 U13877 ( .A(n7965), .B(n8106), .Z(n8223) );
  HS65_LL_IVX9 U13878 ( .A(n3129), .Z(n648) );
  HS65_LL_NAND2X7 U13879 ( .A(n7183), .B(n6476), .Z(n6520) );
  HS65_LL_NAND2X7 U13880 ( .A(n5591), .B(n4883), .Z(n4927) );
  HS65_LL_NOR2X6 U13881 ( .A(n4461), .B(n5532), .Z(n5278) );
  HS65_LL_NOR2X6 U13882 ( .A(n4500), .B(n5554), .Z(n5393) );
  HS65_LL_NOR2X6 U13883 ( .A(n6054), .B(n7124), .Z(n6870) );
  HS65_LL_NOR2X6 U13884 ( .A(n6093), .B(n7146), .Z(n6985) );
  HS65_LL_NOR2X6 U13885 ( .A(n1538), .B(n1544), .Z(n1729) );
  HS65_LL_NOR2X6 U13886 ( .A(n2876), .B(n2969), .Z(n3671) );
  HS65_LL_NOR2X6 U13887 ( .A(n4789), .B(n5555), .Z(n4960) );
  HS65_LL_NOR2X6 U13888 ( .A(n6382), .B(n7147), .Z(n6553) );
  HS65_LL_IVX9 U13889 ( .A(n2913), .Z(n146) );
  HS65_LL_NOR2X6 U13890 ( .A(n3134), .B(n3140), .Z(n3765) );
  HS65_LL_NOR2X6 U13891 ( .A(n7966), .B(n7860), .Z(n8287) );
  HS65_LL_NOR2X6 U13892 ( .A(n3184), .B(n3203), .Z(n3880) );
  HS65_LL_NOR2X6 U13893 ( .A(n2146), .B(n1985), .Z(n1979) );
  HS65_LL_IVX9 U13894 ( .A(n8169), .Z(n123) );
  HS65_LL_IVX9 U13895 ( .A(n8146), .Z(n603) );
  HS65_LL_NOR2X6 U13896 ( .A(n2522), .B(n2361), .Z(n2355) );
  HS65_LL_NOR2X6 U13897 ( .A(n1394), .B(n1233), .Z(n1227) );
  HS65_LL_NOR2X6 U13898 ( .A(n1770), .B(n1609), .Z(n1603) );
  HS65_LL_NOR2X6 U13899 ( .A(n7966), .B(n8082), .Z(n8284) );
  HS65_LL_NOR2X6 U13900 ( .A(n2520), .B(n2289), .Z(n2458) );
  HS65_LL_NOR2X6 U13901 ( .A(n3928), .B(n3096), .Z(n3089) );
  HS65_LL_NOR2X6 U13902 ( .A(n2144), .B(n1913), .Z(n2082) );
  HS65_LL_NOR2X6 U13903 ( .A(n1392), .B(n1161), .Z(n1330) );
  HS65_LL_NOR2X6 U13904 ( .A(n1144), .B(n1180), .Z(n1188) );
  HS65_LL_NOR2X6 U13905 ( .A(n1768), .B(n1537), .Z(n1706) );
  HS65_LL_NOR2X6 U13906 ( .A(n7768), .B(n8527), .Z(n8509) );
  HS65_LL_NOR2X6 U13907 ( .A(n7196), .B(n6475), .Z(n6898) );
  HS65_LL_NOR2X6 U13908 ( .A(n7941), .B(n7942), .Z(n8571) );
  HS65_LL_NOR2X6 U13909 ( .A(n4461), .B(n4747), .Z(n5279) );
  HS65_LL_NOR2X6 U13910 ( .A(n6054), .B(n6327), .Z(n6871) );
  HS65_LL_NOR2X6 U13911 ( .A(n7947), .B(n7769), .Z(n8567) );
  HS65_LL_AOI212X4 U13912 ( .A(n57), .B(n75), .C(n78), .D(n6925), .E(n6057), 
        .Z(n6915) );
  HS65_LL_NAND2X7 U13913 ( .A(n6179), .B(n6516), .Z(n6925) );
  HS65_LL_IVX9 U13914 ( .A(n6926), .Z(n75) );
  HS65_LL_AOI212X4 U13915 ( .A(n579), .B(n601), .C(n612), .D(n8741), .E(n7838), 
        .Z(n8733) );
  HS65_LL_NAND2X7 U13916 ( .A(n7686), .B(n8155), .Z(n8741) );
  HS65_LL_IVX9 U13917 ( .A(n8742), .Z(n601) );
  HS65_LL_NOR2X6 U13918 ( .A(n3972), .B(n3380), .Z(n3374) );
  HS65_LL_NOR2X6 U13919 ( .A(n1163), .B(n1116), .Z(n1335) );
  HS65_LL_NOR2X6 U13920 ( .A(n1915), .B(n1868), .Z(n2087) );
  HS65_LL_NOR2X6 U13921 ( .A(n5591), .B(n5588), .Z(n5319) );
  HS65_LL_NOR2X6 U13922 ( .A(n7183), .B(n7180), .Z(n6911) );
  HS65_LL_NOR2X6 U13923 ( .A(n7208), .B(n7222), .Z(n7026) );
  HS65_LL_NOR2X6 U13924 ( .A(n7971), .B(n7965), .Z(n8232) );
  HS65_LL_NOR2X6 U13925 ( .A(n7948), .B(n8039), .Z(n8590) );
  HS65_LL_NOR2X6 U13926 ( .A(n7847), .B(n7971), .Z(n8288) );
  HS65_LL_NOR2X6 U13927 ( .A(n3952), .B(n3326), .Z(n3320) );
  HS65_LL_NOR2X6 U13928 ( .A(n1539), .B(n1492), .Z(n1711) );
  HS65_LL_NOR2X6 U13929 ( .A(n2291), .B(n2244), .Z(n2463) );
  HS65_LL_NOR2X6 U13930 ( .A(n8033), .B(n8339), .Z(n8600) );
  HS65_LL_NOR2X6 U13931 ( .A(n8039), .B(n8033), .Z(n8534) );
  HS65_LL_NOR2X6 U13932 ( .A(n3731), .B(n3293), .Z(n3309) );
  HS65_LL_NOR2X6 U13933 ( .A(n1487), .B(n1537), .Z(n1648) );
  HS65_LL_NOR2X6 U13934 ( .A(n6348), .B(n6476), .Z(n6893) );
  HS65_LL_NOR2X6 U13935 ( .A(n2831), .B(n3197), .Z(n3787) );
  HS65_LL_NOR2X6 U13936 ( .A(n2239), .B(n2289), .Z(n2400) );
  HS65_LL_NOR2X6 U13937 ( .A(n1863), .B(n1913), .Z(n2024) );
  HS65_LL_NOR2X6 U13938 ( .A(n1111), .B(n1161), .Z(n1272) );
  HS65_LL_NOR2X6 U13939 ( .A(n8123), .B(n8649), .Z(n8292) );
  HS65_LL_NOR2X6 U13940 ( .A(n2497), .B(n2258), .Z(n2319) );
  HS65_LL_AOI212X4 U13941 ( .A(n150), .B(n3597), .C(n154), .D(n174), .E(n4111), 
        .Z(n4108) );
  HS65_LL_CBI4I1X5 U13942 ( .A(n3035), .B(n2918), .C(n3043), .D(n3544), .Z(
        n4111) );
  HS65_LL_NOR2X6 U13943 ( .A(n2121), .B(n1882), .Z(n1943) );
  HS65_LL_NOR2X6 U13944 ( .A(n1369), .B(n1130), .Z(n1191) );
  HS65_LL_NOR2X6 U13945 ( .A(n1745), .B(n1506), .Z(n1567) );
  HS65_LL_NAND2X7 U13946 ( .A(n1909), .B(n2146), .Z(n2052) );
  HS65_LL_NOR2X6 U13947 ( .A(n2969), .B(n3141), .Z(n3766) );
  HS65_LL_NOR2X6 U13948 ( .A(n1522), .B(n1537), .Z(n1734) );
  HS65_LL_NAND2X7 U13949 ( .A(n2285), .B(n2522), .Z(n2428) );
  HS65_LL_NAND2X7 U13950 ( .A(n1157), .B(n1394), .Z(n1300) );
  HS65_LL_NAND2X7 U13951 ( .A(n1533), .B(n1770), .Z(n1676) );
  HS65_LL_NOR2X6 U13952 ( .A(n3116), .B(n3450), .Z(n3445) );
  HS65_LL_NOR2X6 U13953 ( .A(n2274), .B(n2289), .Z(n2486) );
  HS65_LL_NOR2X6 U13954 ( .A(n8556), .B(n8339), .Z(n8334) );
  HS65_LL_NOR2X6 U13955 ( .A(n1146), .B(n1161), .Z(n1358) );
  HS65_LL_NOR2X6 U13956 ( .A(n1898), .B(n1913), .Z(n2110) );
  HS65_LL_NOR2X6 U13957 ( .A(n4733), .B(n5532), .Z(n5298) );
  HS65_LL_NOR2X6 U13958 ( .A(n6329), .B(n7124), .Z(n6890) );
  HS65_LL_NOR2X6 U13959 ( .A(n4591), .B(n4448), .Z(n4917) );
  HS65_LL_NOR2X6 U13960 ( .A(n4608), .B(n4509), .Z(n4970) );
  HS65_LL_NOR2X6 U13961 ( .A(n6201), .B(n6102), .Z(n6563) );
  HS65_LL_NOR2X6 U13962 ( .A(n6184), .B(n6041), .Z(n6510) );
  HS65_LL_NOR2X6 U13963 ( .A(n3141), .B(n3134), .Z(n3724) );
  HS65_LL_NOR2X6 U13964 ( .A(n7836), .B(n8132), .Z(n8716) );
  HS65_LL_NOR2X6 U13965 ( .A(n7875), .B(n8183), .Z(n8806) );
  HS65_LL_NOR2X6 U13966 ( .A(n3342), .B(n2876), .Z(n3155) );
  HS65_LL_NOR2X6 U13967 ( .A(n7180), .B(n7196), .Z(n6860) );
  HS65_LL_NOR2X6 U13968 ( .A(n5588), .B(n5604), .Z(n5268) );
  HS65_LL_NOR2X6 U13969 ( .A(n7943), .B(n8029), .Z(n7954) );
  HS65_LL_NAND2X7 U13970 ( .A(n2240), .B(n2273), .Z(n2287) );
  HS65_LL_NAND2X7 U13971 ( .A(n1488), .B(n1521), .Z(n1535) );
  HS65_LL_NAND2X7 U13972 ( .A(n1864), .B(n1897), .Z(n1911) );
  HS65_LL_NAND2X7 U13973 ( .A(n1112), .B(n1145), .Z(n1159) );
  HS65_LL_NOR2X6 U13974 ( .A(n6054), .B(n7183), .Z(n6921) );
  HS65_LL_NOR2X6 U13975 ( .A(n4461), .B(n5591), .Z(n5329) );
  HS65_LL_NOR2X6 U13976 ( .A(n4500), .B(n5616), .Z(n5444) );
  HS65_LL_NOR2X6 U13977 ( .A(n6093), .B(n7208), .Z(n7036) );
  HS65_LL_NOR4ABX2 U13978 ( .A(n2166), .B(n2167), .C(n2168), .D(n2169), .Z(
        n2133) );
  HS65_LL_OAI222X2 U13979 ( .A(n2144), .B(n1895), .C(n1920), .D(n1897), .E(
        n2069), .F(n1914), .Z(n2169) );
  HS65_LL_NOR3X4 U13980 ( .A(n2032), .B(n1934), .C(n1986), .Z(n2166) );
  HS65_LL_OAI212X5 U13981 ( .A(n2120), .B(n1881), .C(n1898), .D(n1985), .E(
        n2170), .Z(n2168) );
  HS65_LL_NOR4ABX2 U13982 ( .A(n1414), .B(n1415), .C(n1416), .D(n1417), .Z(
        n1381) );
  HS65_LL_OAI222X2 U13983 ( .A(n1392), .B(n1143), .C(n1168), .D(n1145), .E(
        n1317), .F(n1162), .Z(n1417) );
  HS65_LL_NOR3X4 U13984 ( .A(n1280), .B(n1182), .C(n1234), .Z(n1414) );
  HS65_LL_NOR4ABX2 U13985 ( .A(n1322), .B(n1204), .C(n1350), .D(n1333), .Z(
        n1415) );
  HS65_LL_NOR2X6 U13986 ( .A(n8082), .B(n7960), .Z(n8268) );
  HS65_LL_NOR2X6 U13987 ( .A(n4454), .B(n5591), .Z(n5346) );
  HS65_LL_NOR2X6 U13988 ( .A(n4493), .B(n5616), .Z(n5461) );
  HS65_LL_NOR2X6 U13989 ( .A(n6086), .B(n7208), .Z(n7053) );
  HS65_LL_NOR2X6 U13990 ( .A(n6047), .B(n7183), .Z(n6938) );
  HS65_LL_NOR2X6 U13991 ( .A(n1745), .B(n1487), .Z(n1625) );
  HS65_LL_NOR4ABX2 U13992 ( .A(n2542), .B(n2543), .C(n2544), .D(n2545), .Z(
        n2509) );
  HS65_LL_OAI222X2 U13993 ( .A(n2520), .B(n2271), .C(n2296), .D(n2273), .E(
        n2445), .F(n2290), .Z(n2545) );
  HS65_LL_NOR3X4 U13994 ( .A(n2408), .B(n2310), .C(n2362), .Z(n2542) );
  HS65_LL_OAI212X5 U13995 ( .A(n2496), .B(n2257), .C(n2274), .D(n2361), .E(
        n2546), .Z(n2544) );
  HS65_LL_NOR4ABX2 U13996 ( .A(n1790), .B(n1791), .C(n1792), .D(n1793), .Z(
        n1757) );
  HS65_LL_OAI222X2 U13997 ( .A(n1768), .B(n1519), .C(n1544), .D(n1521), .E(
        n1693), .F(n1538), .Z(n1793) );
  HS65_LL_NOR3X4 U13998 ( .A(n1656), .B(n1558), .C(n1610), .Z(n1790) );
  HS65_LL_OAI212X5 U13999 ( .A(n1744), .B(n1505), .C(n1522), .D(n1609), .E(
        n1794), .Z(n1792) );
  HS65_LL_NOR2X6 U14000 ( .A(n2497), .B(n2239), .Z(n2377) );
  HS65_LL_NOR4ABX2 U14001 ( .A(n1175), .B(n1176), .C(n1177), .D(n1178), .Z(
        n1137) );
  HS65_LL_OAI212X5 U14002 ( .A(n1112), .B(n1179), .C(n1162), .D(n1180), .E(
        n1181), .Z(n1178) );
  HS65_LL_NAND3AX6 U14003 ( .A(n1182), .B(n1183), .C(n1184), .Z(n1177) );
  HS65_LL_NOR3AX2 U14004 ( .A(n1190), .B(n1191), .C(n1192), .Z(n1175) );
  HS65_LL_NOR4ABX2 U14005 ( .A(n1927), .B(n1928), .C(n1929), .D(n1930), .Z(
        n1889) );
  HS65_LL_OAI212X5 U14006 ( .A(n1864), .B(n1931), .C(n1914), .D(n1932), .E(
        n1933), .Z(n1930) );
  HS65_LL_NAND3AX6 U14007 ( .A(n1934), .B(n1935), .C(n1936), .Z(n1929) );
  HS65_LL_NOR3AX2 U14008 ( .A(n1942), .B(n1943), .C(n1944), .Z(n1927) );
  HS65_LL_NOR2X6 U14009 ( .A(n1369), .B(n1111), .Z(n1249) );
  HS65_LL_NOR2X6 U14010 ( .A(n2121), .B(n1863), .Z(n2001) );
  HS65_LL_NOR4ABX2 U14011 ( .A(n2303), .B(n2304), .C(n2305), .D(n2306), .Z(
        n2265) );
  HS65_LL_NAND3AX6 U14012 ( .A(n2310), .B(n2311), .C(n2312), .Z(n2305) );
  HS65_LL_OAI212X5 U14013 ( .A(n2240), .B(n2307), .C(n2290), .D(n2308), .E(
        n2309), .Z(n2306) );
  HS65_LL_NOR3AX2 U14014 ( .A(n2318), .B(n2319), .C(n2320), .Z(n2303) );
  HS65_LL_NOR4ABX2 U14015 ( .A(n1551), .B(n1552), .C(n1553), .D(n1554), .Z(
        n1513) );
  HS65_LL_NAND3AX6 U14016 ( .A(n1558), .B(n1559), .C(n1560), .Z(n1553) );
  HS65_LL_NOR4ABX2 U14017 ( .A(n1562), .B(n1563), .C(n1564), .D(n1565), .Z(
        n1552) );
  HS65_LL_OAI212X5 U14018 ( .A(n1488), .B(n1555), .C(n1538), .D(n1556), .E(
        n1557), .Z(n1554) );
  HS65_LL_NOR2X6 U14019 ( .A(n7960), .B(n8106), .Z(n8291) );
  HS65_LL_NOR2X6 U14020 ( .A(n3972), .B(n2993), .Z(n3847) );
  HS65_LL_NOR2X6 U14021 ( .A(n3952), .B(n2968), .Z(n3732) );
  HS65_LL_NOR2X6 U14022 ( .A(n6348), .B(n6055), .Z(n6900) );
  HS65_LL_NOR2X6 U14023 ( .A(n4732), .B(n4462), .Z(n5308) );
  HS65_LL_NOR2X6 U14024 ( .A(n4794), .B(n4501), .Z(n5423) );
  HS65_LL_NOR2X6 U14025 ( .A(n6387), .B(n6094), .Z(n7015) );
  HS65_LL_CBI4I1X5 U14026 ( .A(n1199), .B(n1180), .C(n1116), .D(n1303), .Z(
        n1302) );
  HS65_LL_CBI4I1X5 U14027 ( .A(n1951), .B(n1932), .C(n1868), .D(n2055), .Z(
        n2054) );
  HS65_LL_NOR2X6 U14028 ( .A(n7821), .B(n7631), .Z(n7792) );
  HS65_LL_NOR2X6 U14029 ( .A(n7919), .B(n7651), .Z(n7891) );
  HS65_LL_NOR2X6 U14030 ( .A(n4789), .B(n4508), .Z(n5397) );
  HS65_LL_NOR2X6 U14031 ( .A(n6382), .B(n6101), .Z(n6989) );
  HS65_LL_NOR2X6 U14032 ( .A(n4727), .B(n4447), .Z(n5282) );
  HS65_LL_NOR2X6 U14033 ( .A(n6343), .B(n6040), .Z(n6874) );
  HS65_LL_NOR2X6 U14034 ( .A(n4643), .B(n4654), .Z(n5165) );
  HS65_LL_NOR2X6 U14035 ( .A(n6236), .B(n6247), .Z(n6757) );
  HS65_LL_NOR2X6 U14036 ( .A(n1985), .B(n1909), .Z(n2032) );
  HS65_LL_NOR2X6 U14037 ( .A(n1233), .B(n1157), .Z(n1280) );
  HS65_LL_NOR2X6 U14038 ( .A(n7147), .B(n6203), .Z(n6538) );
  HS65_LL_NOR2X6 U14039 ( .A(n7125), .B(n6186), .Z(n6485) );
  HS65_LL_NOR2X6 U14040 ( .A(n5533), .B(n4593), .Z(n4892) );
  HS65_LL_NOR2X6 U14041 ( .A(n5555), .B(n4610), .Z(n4945) );
  HS65_LL_CBI4I1X5 U14042 ( .A(n2327), .B(n2308), .C(n2244), .D(n2431), .Z(
        n2430) );
  HS65_LL_CBI4I1X5 U14043 ( .A(n1575), .B(n1556), .C(n1492), .D(n1679), .Z(
        n1678) );
  HS65_LL_NOR2X6 U14044 ( .A(n2361), .B(n2285), .Z(n2408) );
  HS65_LL_NOR2X6 U14045 ( .A(n1609), .B(n1533), .Z(n1656) );
  HS65_LL_NOR4ABX2 U14046 ( .A(n1735), .B(n1736), .C(n1737), .D(n1738), .Z(
        n1582) );
  HS65_LL_NOR3X4 U14047 ( .A(n1747), .B(n1748), .C(n1749), .Z(n1736) );
  HS65_LL_NAND4ABX3 U14048 ( .A(n1739), .B(n1496), .C(n1740), .D(n1741), .Z(
        n1738) );
  HS65_LL_OAI212X5 U14049 ( .A(n1742), .B(n1743), .C(n1744), .D(n1745), .E(
        n1746), .Z(n1737) );
  HS65_LL_NOR4ABX2 U14050 ( .A(n2487), .B(n2488), .C(n2489), .D(n2490), .Z(
        n2334) );
  HS65_LL_NOR3X4 U14051 ( .A(n2499), .B(n2500), .C(n2501), .Z(n2488) );
  HS65_LL_OAI212X5 U14052 ( .A(n2494), .B(n2495), .C(n2496), .D(n2497), .E(
        n2498), .Z(n2489) );
  HS65_LL_NAND4ABX3 U14053 ( .A(n2491), .B(n2248), .C(n2492), .D(n2493), .Z(
        n2490) );
  HS65_LL_NOR4ABX2 U14054 ( .A(n2111), .B(n2112), .C(n2113), .D(n2114), .Z(
        n1958) );
  HS65_LL_NOR3X4 U14055 ( .A(n2123), .B(n2124), .C(n2125), .Z(n2112) );
  HS65_LL_OAI212X5 U14056 ( .A(n2118), .B(n2119), .C(n2120), .D(n2121), .E(
        n2122), .Z(n2113) );
  HS65_LL_NAND4ABX3 U14057 ( .A(n2115), .B(n1872), .C(n2116), .D(n2117), .Z(
        n2114) );
  HS65_LL_NOR4ABX2 U14058 ( .A(n1359), .B(n1360), .C(n1361), .D(n1362), .Z(
        n1206) );
  HS65_LL_NOR3X4 U14059 ( .A(n1371), .B(n1372), .C(n1373), .Z(n1360) );
  HS65_LL_NAND4ABX3 U14060 ( .A(n1363), .B(n1120), .C(n1364), .D(n1365), .Z(
        n1362) );
  HS65_LL_OAI212X5 U14061 ( .A(n1366), .B(n1367), .C(n1368), .D(n1369), .E(
        n1370), .Z(n1361) );
  HS65_LL_NOR2X6 U14062 ( .A(n1770), .B(n1520), .Z(n1696) );
  HS65_LL_NOR2X6 U14063 ( .A(n2522), .B(n2272), .Z(n2448) );
  HS65_LL_NOR2X6 U14064 ( .A(n1394), .B(n1144), .Z(n1320) );
  HS65_LL_NOR2X6 U14065 ( .A(n2146), .B(n1896), .Z(n2072) );
  HS65_LL_NOR2X6 U14066 ( .A(n2276), .B(n2520), .Z(n2330) );
  HS65_LL_NOR2X6 U14067 ( .A(n1900), .B(n2144), .Z(n1954) );
  HS65_LL_NOR2X6 U14068 ( .A(n1148), .B(n1392), .Z(n1202) );
  HS65_LL_NAND2X7 U14069 ( .A(n8776), .B(n8449), .Z(n8756) );
  HS65_LL_NAND2X7 U14070 ( .A(n8686), .B(n8397), .Z(n8666) );
  HS65_LL_NOR2X6 U14071 ( .A(n1524), .B(n1768), .Z(n1578) );
  HS65_LL_NOR2X6 U14072 ( .A(n3396), .B(n2831), .Z(n3400) );
  HS65_LL_NOR2X6 U14073 ( .A(n2830), .B(n3204), .Z(n3802) );
  HS65_LL_NOR2X6 U14074 ( .A(n2307), .B(n2333), .Z(n2442) );
  HS65_LL_NOR2X6 U14075 ( .A(n1555), .B(n1581), .Z(n1690) );
  HS65_LL_NOR2X6 U14076 ( .A(n1179), .B(n1205), .Z(n1314) );
  HS65_LL_NOR2X6 U14077 ( .A(n1931), .B(n1957), .Z(n2066) );
  HS65_LL_NOR2X6 U14078 ( .A(n1145), .B(n1180), .Z(n1275) );
  HS65_LL_NOR2X6 U14079 ( .A(n1897), .B(n1932), .Z(n2027) );
  HS65_LL_NOR2X6 U14080 ( .A(n2859), .B(n3926), .Z(n3064) );
  HS65_LL_NOR2X6 U14081 ( .A(n2997), .B(n3970), .Z(n3409) );
  HS65_LL_NOR2X6 U14082 ( .A(n7949), .B(n8028), .Z(n8333) );
  HS65_LL_NOR2X6 U14083 ( .A(n2273), .B(n2308), .Z(n2403) );
  HS65_LL_NOR2X6 U14084 ( .A(n3342), .B(n2883), .Z(n3346) );
  HS65_LL_NOR2X6 U14085 ( .A(n1521), .B(n1556), .Z(n1651) );
  HS65_LL_NOR2X6 U14086 ( .A(n8123), .B(n7993), .Z(n8307) );
  HS65_LL_NOR2X6 U14087 ( .A(n7750), .B(n8082), .Z(n7991) );
  HS65_LL_NOR2X6 U14088 ( .A(n7947), .B(n8339), .Z(n8059) );
  HS65_LL_NOR2X6 U14089 ( .A(n1868), .B(n1920), .Z(n2092) );
  HS65_LL_NOR2X6 U14090 ( .A(n1116), .B(n1168), .Z(n1340) );
  HS65_LL_NOR4ABX2 U14091 ( .A(n2135), .B(n2136), .C(n2137), .D(n2138), .Z(
        n1878) );
  HS65_LL_CBI4I1X5 U14092 ( .A(n1881), .B(n1957), .C(n1898), .D(n1977), .Z(
        n2137) );
  HS65_LL_CBI4I1X5 U14093 ( .A(n2056), .B(n1921), .C(n1868), .D(n2139), .Z(
        n2138) );
  HS65_LL_NOR4ABX2 U14094 ( .A(n2022), .B(n2061), .C(n2082), .D(n2105), .Z(
        n2135) );
  HS65_LL_NOR4ABX2 U14095 ( .A(n1383), .B(n1384), .C(n1385), .D(n1386), .Z(
        n1126) );
  HS65_LL_CBI4I1X5 U14096 ( .A(n1129), .B(n1205), .C(n1146), .D(n1225), .Z(
        n1385) );
  HS65_LL_CBI4I1X5 U14097 ( .A(n1304), .B(n1169), .C(n1116), .D(n1387), .Z(
        n1386) );
  HS65_LL_NOR4ABX2 U14098 ( .A(n1270), .B(n1309), .C(n1330), .D(n1353), .Z(
        n1383) );
  HS65_LL_NOR4ABX2 U14099 ( .A(n2511), .B(n2512), .C(n2513), .D(n2514), .Z(
        n2254) );
  HS65_LL_CBI4I1X5 U14100 ( .A(n2257), .B(n2333), .C(n2274), .D(n2353), .Z(
        n2513) );
  HS65_LL_CBI4I1X5 U14101 ( .A(n2432), .B(n2297), .C(n2244), .D(n2515), .Z(
        n2514) );
  HS65_LL_NOR4ABX2 U14102 ( .A(n2398), .B(n2437), .C(n2458), .D(n2481), .Z(
        n2511) );
  HS65_LL_NOR4ABX2 U14103 ( .A(n1759), .B(n1760), .C(n1761), .D(n1762), .Z(
        n1502) );
  HS65_LL_CBI4I1X5 U14104 ( .A(n1505), .B(n1581), .C(n1522), .D(n1601), .Z(
        n1761) );
  HS65_LL_CBI4I1X5 U14105 ( .A(n1680), .B(n1545), .C(n1492), .D(n1763), .Z(
        n1762) );
  HS65_LL_NOR4ABX2 U14106 ( .A(n1646), .B(n1685), .C(n1706), .D(n1729), .Z(
        n1759) );
  HS65_LL_NOR2X6 U14107 ( .A(n1492), .B(n1544), .Z(n1716) );
  HS65_LL_NOR2X6 U14108 ( .A(n2244), .B(n2296), .Z(n2468) );
  HS65_LL_NOR2X6 U14109 ( .A(n1544), .B(n1532), .Z(n1639) );
  HS65_LL_NOR2X6 U14110 ( .A(n2361), .B(n2297), .Z(n2345) );
  HS65_LL_NAND2X7 U14111 ( .A(n1745), .B(n1493), .Z(n1661) );
  HS65_LL_NOR2X6 U14112 ( .A(n3475), .B(n2938), .Z(n3513) );
  HS65_LL_NOR2X6 U14113 ( .A(n1985), .B(n1921), .Z(n1969) );
  HS65_LL_NOR2X6 U14114 ( .A(n1233), .B(n1169), .Z(n1217) );
  HS65_LL_NOR2X6 U14115 ( .A(n2296), .B(n2284), .Z(n2391) );
  HS65_LL_NOR2X6 U14116 ( .A(n1920), .B(n1908), .Z(n2015) );
  HS65_LL_NOR2X6 U14117 ( .A(n1168), .B(n1156), .Z(n1263) );
  HS65_LL_NAND2X7 U14118 ( .A(n2497), .B(n2245), .Z(n2413) );
  HS65_LL_NAND2X7 U14119 ( .A(n2121), .B(n1869), .Z(n2037) );
  HS65_LL_NAND2X7 U14120 ( .A(n1369), .B(n1117), .Z(n1285) );
  HS65_LL_NOR2X6 U14121 ( .A(n7965), .B(n7860), .Z(n8248) );
  HS65_LL_NOR2X6 U14122 ( .A(n1494), .B(n1524), .Z(n1614) );
  HS65_LL_NOR2X6 U14123 ( .A(n2246), .B(n2276), .Z(n2366) );
  HS65_LL_NOR2X6 U14124 ( .A(n1118), .B(n1148), .Z(n1238) );
  HS65_LL_NOR2X6 U14125 ( .A(n1870), .B(n1900), .Z(n1990) );
  HS65_LL_NOR2X6 U14126 ( .A(n2882), .B(n3692), .Z(n3675) );
  HS65_LL_NOR2X6 U14127 ( .A(n8033), .B(n7942), .Z(n8550) );
  HS65_LL_NOR2X6 U14128 ( .A(n2829), .B(n3412), .Z(n3826) );
  HS65_LL_NOR2X6 U14129 ( .A(n8173), .B(n7875), .Z(n8802) );
  HS65_LL_NOR2X6 U14130 ( .A(n8150), .B(n7836), .Z(n8712) );
  HS65_LL_NAND2X7 U14131 ( .A(n1537), .B(n1493), .Z(n1594) );
  HS65_LL_NOR2X6 U14132 ( .A(n2071), .B(n1920), .Z(n2073) );
  HS65_LL_NOR2X6 U14133 ( .A(n1319), .B(n1168), .Z(n1321) );
  HS65_LL_NAND2X7 U14134 ( .A(n2289), .B(n2245), .Z(n2346) );
  HS65_LL_NAND2X7 U14135 ( .A(n1161), .B(n1117), .Z(n1218) );
  HS65_LL_NAND2X7 U14136 ( .A(n1913), .B(n1869), .Z(n1970) );
  HS65_LL_NOR2X6 U14137 ( .A(n2981), .B(n3141), .Z(n3349) );
  HS65_LL_NOR2X6 U14138 ( .A(n6260), .B(n6076), .Z(n6657) );
  HS65_LL_NOR2X6 U14139 ( .A(n4667), .B(n4483), .Z(n5064) );
  HS65_LL_NOR2X6 U14140 ( .A(n4994), .B(n4501), .Z(n5417) );
  HS65_LL_NOR2X6 U14141 ( .A(n6587), .B(n6094), .Z(n7009) );
  HS65_LL_NOR2X6 U14142 ( .A(n4882), .B(n4462), .Z(n5302) );
  HS65_LL_NOR2X6 U14143 ( .A(n6475), .B(n6055), .Z(n6894) );
  HS65_LL_NOR2X6 U14144 ( .A(n8302), .B(n7859), .Z(n8297) );
  HS65_LL_NOR2X6 U14145 ( .A(n2447), .B(n2296), .Z(n2449) );
  HS65_LL_NOR2X6 U14146 ( .A(n8034), .B(n7769), .Z(n8589) );
  HS65_LL_NOR2X6 U14147 ( .A(n1695), .B(n1544), .Z(n1697) );
  HS65_LL_NAND2X7 U14148 ( .A(n2119), .B(n1898), .Z(n1989) );
  HS65_LL_NOR2X6 U14149 ( .A(n1743), .B(n1745), .Z(n1663) );
  HS65_LL_NOR2X6 U14150 ( .A(n8357), .B(n7948), .Z(n8599) );
  HS65_LL_NOR2AX3 U14151 ( .A(n6182), .B(n6184), .Z(n6852) );
  HS65_LL_NOR2AX3 U14152 ( .A(n4589), .B(n4591), .Z(n5260) );
  HS65_LL_NOR2AX3 U14153 ( .A(n4606), .B(n4608), .Z(n5375) );
  HS65_LL_NOR2AX3 U14154 ( .A(n6199), .B(n6201), .Z(n6967) );
  HS65_LL_NOR2X6 U14155 ( .A(n2495), .B(n2497), .Z(n2415) );
  HS65_LL_NOR2X6 U14156 ( .A(n2119), .B(n2121), .Z(n2039) );
  HS65_LL_NOR2X6 U14157 ( .A(n1367), .B(n1369), .Z(n1287) );
  HS65_LL_NOR2X6 U14158 ( .A(n1861), .B(n1957), .Z(n2049) );
  HS65_LL_NAND2X7 U14159 ( .A(n2495), .B(n2274), .Z(n2365) );
  HS65_LL_NAND2X7 U14160 ( .A(n1367), .B(n1146), .Z(n1237) );
  HS65_LL_NAND2X7 U14161 ( .A(n1743), .B(n1522), .Z(n1613) );
  HS65_LL_NOR2X6 U14162 ( .A(n2237), .B(n2333), .Z(n2425) );
  HS65_LL_NOR2X6 U14163 ( .A(n1109), .B(n1205), .Z(n1297) );
  HS65_LL_NOR2X6 U14164 ( .A(n1485), .B(n1581), .Z(n1673) );
  HS65_LL_NOR2X6 U14165 ( .A(n3846), .B(n3203), .Z(n3848) );
  HS65_LL_NOR2X6 U14166 ( .A(n1117), .B(n1168), .Z(n1336) );
  HS65_LL_NOR2X6 U14167 ( .A(n1869), .B(n1920), .Z(n2088) );
  HS65_LL_NAND4ABX3 U14168 ( .A(n7681), .B(n575), .C(n7682), .D(n7683), .Z(
        n7629) );
  HS65_LL_NOR3AX2 U14169 ( .A(n7688), .B(n7689), .C(n7690), .Z(n7682) );
  HS65_LL_AOI212X4 U14170 ( .A(n614), .B(n7684), .C(n587), .D(n617), .E(n7685), 
        .Z(n7683) );
  HS65_LL_MX41X7 U14171 ( .D0(n591), .S0(n612), .D1(n585), .S1(n609), .D2(n615), .S2(n578), .D3(n605), .S3(n7699), .Z(n7681) );
  HS65_LL_NAND4ABX3 U14172 ( .A(n7719), .B(n95), .C(n7720), .D(n7721), .Z(
        n7649) );
  HS65_LL_NOR3AX2 U14173 ( .A(n7726), .B(n7727), .C(n7728), .Z(n7720) );
  HS65_LL_AOI212X4 U14174 ( .A(n134), .B(n7722), .C(n107), .D(n137), .E(n7723), 
        .Z(n7721) );
  HS65_LL_MX41X7 U14175 ( .D0(n111), .S0(n132), .D1(n105), .S1(n129), .D2(n135), .S2(n98), .D3(n125), .S3(n7737), .Z(n7719) );
  HS65_LL_NOR2X6 U14176 ( .A(n7768), .B(n8357), .Z(n8060) );
  HS65_LL_NOR2X6 U14177 ( .A(n7622), .B(n8150), .Z(n7672) );
  HS65_LL_NOR2X6 U14178 ( .A(n2881), .B(n3299), .Z(n3711) );
  HS65_LL_NOR2X6 U14179 ( .A(n2245), .B(n2296), .Z(n2464) );
  HS65_LL_NOR2X6 U14180 ( .A(n7630), .B(n7676), .Z(n7789) );
  HS65_LL_NOR2X6 U14181 ( .A(n1493), .B(n1544), .Z(n1712) );
  HS65_LL_NOR2X6 U14182 ( .A(n2938), .B(n2926), .Z(n3419) );
  HS65_LL_NOR2X6 U14183 ( .A(n8067), .B(n8207), .Z(n7746) );
  HS65_LL_NOR2X6 U14184 ( .A(n7850), .B(n8106), .Z(n8270) );
  HS65_LL_NOR2X6 U14185 ( .A(n2307), .B(n2257), .Z(n2360) );
  HS65_LL_NOR2X6 U14186 ( .A(n1555), .B(n1505), .Z(n1608) );
  HS65_LL_NOR2X6 U14187 ( .A(n1931), .B(n1881), .Z(n1984) );
  HS65_LL_NOR2X6 U14188 ( .A(n1179), .B(n1129), .Z(n1232) );
  HS65_LL_NOR2X6 U14189 ( .A(n2882), .B(n3141), .Z(n3687) );
  HS65_LL_IVX9 U14190 ( .A(n8776), .Z(n113) );
  HS65_LL_NOR2X6 U14191 ( .A(n2836), .B(n3203), .Z(n3867) );
  HS65_LL_NOR2X6 U14192 ( .A(n2837), .B(n3203), .Z(n3863) );
  HS65_LL_NOR2X6 U14193 ( .A(n2071), .B(n1951), .Z(n1968) );
  HS65_LL_NOR2X6 U14194 ( .A(n1985), .B(n1951), .Z(n1992) );
  HS65_LL_NOR2X6 U14195 ( .A(n1319), .B(n1199), .Z(n1216) );
  HS65_LL_NOR2X6 U14196 ( .A(n1233), .B(n1199), .Z(n1240) );
  HS65_LL_NOR2X6 U14197 ( .A(n1533), .B(n1581), .Z(n1495) );
  HS65_LL_NOR2X6 U14198 ( .A(n2285), .B(n2333), .Z(n2247) );
  HS65_LL_NOR2X6 U14199 ( .A(n1157), .B(n1205), .Z(n1119) );
  HS65_LL_NOR2X6 U14200 ( .A(n1909), .B(n1957), .Z(n1871) );
  HS65_LL_NOR2X6 U14201 ( .A(n1881), .B(n1863), .Z(n1941) );
  HS65_LL_NOR2X6 U14202 ( .A(n1864), .B(n1861), .Z(n2065) );
  HS65_LL_NOR2X6 U14203 ( .A(n1556), .B(n1581), .Z(n1568) );
  HS65_LL_NOR2X6 U14204 ( .A(n2308), .B(n2333), .Z(n2320) );
  HS65_LL_NOR2X6 U14205 ( .A(n1180), .B(n1205), .Z(n1192) );
  HS65_LL_NOR2X6 U14206 ( .A(n1932), .B(n1957), .Z(n1944) );
  HS65_LL_CBI4I1X5 U14207 ( .A(n3293), .B(n3158), .C(n2888), .D(n3716), .Z(
        n3715) );
  HS65_LL_NOR4ABX2 U14208 ( .A(n7197), .B(n7198), .C(n7199), .D(n7200), .Z(
        n7113) );
  HS65_LL_OAI222X2 U14209 ( .A(n6186), .B(n7196), .C(n7124), .D(n6515), .E(
        n6857), .F(n6329), .Z(n7200) );
  HS65_LL_NOR3X4 U14210 ( .A(n6337), .B(n6887), .C(n6931), .Z(n7197) );
  HS65_LL_OAI212X5 U14211 ( .A(n6926), .B(n6041), .C(n6516), .D(n6476), .E(
        n7201), .Z(n7199) );
  HS65_LL_NOR2X6 U14212 ( .A(n3731), .B(n3140), .Z(n3733) );
  HS65_LL_NOR2X6 U14213 ( .A(n2272), .B(n2258), .Z(n2375) );
  HS65_LL_NOR2X6 U14214 ( .A(n8630), .B(n7767), .Z(n8605) );
  HS65_LL_NOR2X6 U14215 ( .A(n1112), .B(n1109), .Z(n1313) );
  HS65_LL_NOR2X6 U14216 ( .A(n1488), .B(n1485), .Z(n1689) );
  HS65_LL_NOR2X6 U14217 ( .A(n2240), .B(n2237), .Z(n2441) );
  HS65_LL_NOR2X6 U14218 ( .A(n2447), .B(n2327), .Z(n2344) );
  HS65_LL_NOR2X6 U14219 ( .A(n2361), .B(n2327), .Z(n2368) );
  HS65_LL_NOR2X6 U14220 ( .A(n1129), .B(n1111), .Z(n1189) );
  HS65_LL_NOR2X6 U14221 ( .A(n2257), .B(n2239), .Z(n2317) );
  HS65_LL_NOR2X6 U14222 ( .A(n1505), .B(n1487), .Z(n1565) );
  HS65_LL_NOR2X6 U14223 ( .A(n1896), .B(n1882), .Z(n1999) );
  HS65_LL_NOR2X6 U14224 ( .A(n1144), .B(n1130), .Z(n1247) );
  HS65_LL_NAND2X7 U14225 ( .A(n5588), .B(n4461), .Z(n5315) );
  HS65_LL_NAND2X7 U14226 ( .A(n7180), .B(n6054), .Z(n6907) );
  HS65_LL_NOR4ABX2 U14227 ( .A(n4014), .B(n4015), .C(n4016), .D(n4017), .Z(
        n3937) );
  HS65_LL_OAI222X2 U14228 ( .A(n3950), .B(n2981), .C(n3140), .D(n2969), .E(
        n3343), .F(n3134), .Z(n4017) );
  HS65_LL_NOR3X4 U14229 ( .A(n3680), .B(n3160), .C(n3327), .Z(n4014) );
  HS65_LL_OAI212X5 U14230 ( .A(n3693), .B(n2875), .C(n2970), .D(n3326), .E(
        n4018), .Z(n4016) );
  HS65_LL_NOR2X6 U14231 ( .A(n7769), .B(n8369), .Z(n8535) );
  HS65_LL_NOR2X6 U14232 ( .A(n1609), .B(n1575), .Z(n1616) );
  HS65_LL_NOR2X6 U14233 ( .A(n1695), .B(n1575), .Z(n1592) );
  HS65_LL_NOR2X6 U14234 ( .A(n1520), .B(n1506), .Z(n1623) );
  HS65_LL_NOR2X6 U14235 ( .A(n3380), .B(n3406), .Z(n3387) );
  HS65_LL_NOR2X6 U14236 ( .A(n8039), .B(n7951), .Z(n8036) );
  HS65_LL_NOR2X6 U14237 ( .A(n2993), .B(n2846), .Z(n3398) );
  HS65_LL_NOR2X6 U14238 ( .A(n2855), .B(n3112), .Z(n3117) );
  HS65_LL_NOR2X6 U14239 ( .A(n2845), .B(n2831), .Z(n3179) );
  HS65_LL_NOR2X6 U14240 ( .A(n1110), .B(n1199), .Z(n1262) );
  HS65_LL_NOR2X6 U14241 ( .A(n1862), .B(n1951), .Z(n2014) );
  HS65_LL_NAND4ABX3 U14242 ( .A(n8624), .B(n8625), .C(n8626), .D(n8627), .Z(
        n7773) );
  HS65_LL_OAI222X2 U14243 ( .A(n8363), .B(n8540), .C(n8556), .D(n7949), .E(
        n7769), .F(n8510), .Z(n8624) );
  HS65_LL_NOR3AX2 U14244 ( .A(n8501), .B(n8552), .C(n8594), .Z(n8626) );
  HS65_LL_NAND4ABX3 U14245 ( .A(n8061), .B(n8338), .C(n8607), .D(n8568), .Z(
        n8625) );
  HS65_LL_NOR2X6 U14246 ( .A(n8649), .B(n7749), .Z(n8218) );
  HS65_LL_NOR2X6 U14247 ( .A(n2447), .B(n2520), .Z(n2376) );
  HS65_LL_NOR2X6 U14248 ( .A(n8117), .B(n8254), .Z(n8090) );
  HS65_LL_NOR2X6 U14249 ( .A(n2258), .B(n2447), .Z(n2462) );
  HS65_LL_IVX9 U14250 ( .A(n8540), .Z(n322) );
  HS65_LL_NOR2X6 U14251 ( .A(n2238), .B(n2327), .Z(n2390) );
  HS65_LL_NOR2X6 U14252 ( .A(n8363), .B(n8556), .Z(n8322) );
  HS65_LL_NOR2X6 U14253 ( .A(n1882), .B(n2071), .Z(n2086) );
  HS65_LL_NOR2X6 U14254 ( .A(n1130), .B(n1319), .Z(n1334) );
  HS65_LL_NOR2X6 U14255 ( .A(n2071), .B(n2144), .Z(n2000) );
  HS65_LL_NOR2X6 U14256 ( .A(n1319), .B(n1392), .Z(n1248) );
  HS65_LL_NOR2X6 U14257 ( .A(n2889), .B(n3157), .Z(n3751) );
  HS65_LL_NOR2X6 U14258 ( .A(n3982), .B(n3042), .Z(n3543) );
  HS65_LL_NOR2X6 U14259 ( .A(n1486), .B(n1575), .Z(n1638) );
  HS65_LL_NOR2X6 U14260 ( .A(n2968), .B(n2876), .Z(n3344) );
  HS65_LL_NAND4ABX3 U14261 ( .A(n8652), .B(n8653), .C(n8654), .D(n8655), .Z(
        n7755) );
  HS65_LL_OAI222X2 U14262 ( .A(n8117), .B(n8238), .C(n8254), .D(n7848), .E(
        n7751), .F(n8207), .Z(n8652) );
  HS65_LL_NAND4ABX3 U14263 ( .A(n7990), .B(n8225), .C(n8103), .D(n8266), .Z(
        n8653) );
  HS65_LL_NOR3AX2 U14264 ( .A(n8198), .B(n8251), .C(n8292), .Z(n8654) );
  HS65_LL_IVX9 U14265 ( .A(n7749), .Z(n365) );
  HS65_LL_NOR2X6 U14266 ( .A(n1506), .B(n1695), .Z(n1710) );
  HS65_LL_NOR2X6 U14267 ( .A(n2889), .B(n3140), .Z(n3748) );
  HS65_LL_NOR2X6 U14268 ( .A(n2888), .B(n3140), .Z(n3752) );
  HS65_LL_NOR2X6 U14269 ( .A(n1695), .B(n1768), .Z(n1624) );
  HS65_LL_NOR2X6 U14270 ( .A(n2875), .B(n2883), .Z(n3153) );
  HS65_LL_NOR2X6 U14271 ( .A(n3096), .B(n3061), .Z(n3104) );
  HS65_LL_NOR2X6 U14272 ( .A(n1555), .B(n1695), .Z(n1691) );
  HS65_LL_NOR2X6 U14273 ( .A(n2307), .B(n2447), .Z(n2443) );
  HS65_LL_NOR2X6 U14274 ( .A(n2308), .B(n2276), .Z(n2424) );
  HS65_LL_NOR2X6 U14275 ( .A(n1556), .B(n1524), .Z(n1672) );
  HS65_LL_NOR2X6 U14276 ( .A(n1180), .B(n1148), .Z(n1296) );
  HS65_LL_NOR2X6 U14277 ( .A(n1932), .B(n1900), .Z(n2048) );
  HS65_LL_NOR2X6 U14278 ( .A(n1179), .B(n1319), .Z(n1315) );
  HS65_LL_NOR2X6 U14279 ( .A(n1931), .B(n2071), .Z(n2067) );
  HS65_LL_NOR2X6 U14280 ( .A(n8556), .B(n8630), .Z(n8361) );
  HS65_LL_NOR2X6 U14281 ( .A(n2940), .B(n3095), .Z(n2952) );
  HS65_LL_NOR2X6 U14282 ( .A(n2846), .B(n3846), .Z(n3861) );
  HS65_LL_NOR2X6 U14283 ( .A(n7860), .B(n8238), .Z(n8275) );
  HS65_LL_NOR2X6 U14284 ( .A(n3846), .B(n3970), .Z(n3399) );
  HS65_LL_NOR2X6 U14285 ( .A(n3491), .B(n3926), .Z(n3118) );
  HS65_LL_NOR2X6 U14286 ( .A(n3135), .B(n2888), .Z(n3747) );
  HS65_LL_NOR2X6 U14287 ( .A(n7859), .B(n7980), .Z(n8274) );
  HS65_LL_CBI4I1X5 U14288 ( .A(n1488), .B(n1524), .C(n1575), .D(n1654), .Z(
        n1808) );
  HS65_LL_CBI4I1X5 U14289 ( .A(n2240), .B(n2276), .C(n2327), .D(n2406), .Z(
        n2560) );
  HS65_LL_CBI4I1X5 U14290 ( .A(n1112), .B(n1148), .C(n1199), .D(n1278), .Z(
        n1432) );
  HS65_LL_CBI4I1X5 U14291 ( .A(n1864), .B(n1900), .C(n1951), .D(n2030), .Z(
        n2184) );
  HS65_LL_NOR2X6 U14292 ( .A(n7941), .B(n8048), .Z(n8575) );
  HS65_LL_NOR2X6 U14293 ( .A(n7846), .B(n7961), .Z(n8273) );
  HS65_LL_NOR2X6 U14294 ( .A(n1862), .B(n2119), .Z(n2028) );
  HS65_LL_NOR2X6 U14295 ( .A(n1869), .B(n2119), .Z(n2115) );
  HS65_LL_NOR2X6 U14296 ( .A(n2876), .B(n3731), .Z(n3746) );
  HS65_LL_NOR2X6 U14297 ( .A(n8146), .B(n8686), .Z(n8152) );
  HS65_LL_NOR2X6 U14298 ( .A(n8169), .B(n8776), .Z(n8175) );
  HS65_LL_IVX9 U14299 ( .A(n2940), .Z(n190) );
  HS65_LL_NOR2X6 U14300 ( .A(n2146), .B(n1881), .Z(n1980) );
  HS65_LL_NOR2X6 U14301 ( .A(n4499), .B(n5380), .Z(n5433) );
  HS65_LL_NOR2X6 U14302 ( .A(n6092), .B(n6972), .Z(n7025) );
  HS65_LL_NOR2X6 U14303 ( .A(n3731), .B(n3950), .Z(n3345) );
  HS65_LL_IVX9 U14304 ( .A(n2274), .Z(n895) );
  HS65_LL_IVX9 U14305 ( .A(n1146), .Z(n854) );
  HS65_LL_IVX9 U14306 ( .A(n1898), .Z(n772) );
  HS65_LL_IVX9 U14307 ( .A(n8207), .Z(n373) );
  HS65_LL_NOR2X6 U14308 ( .A(n1110), .B(n1367), .Z(n1276) );
  HS65_LL_NOR2X6 U14309 ( .A(n2238), .B(n2495), .Z(n2404) );
  HS65_LL_NOR2X6 U14310 ( .A(n1486), .B(n1743), .Z(n1652) );
  HS65_LL_NOR2X6 U14311 ( .A(n2245), .B(n2495), .Z(n2491) );
  HS65_LL_NOR2X6 U14312 ( .A(n1117), .B(n1367), .Z(n1363) );
  HS65_LL_NOR2X6 U14313 ( .A(n1493), .B(n1743), .Z(n1739) );
  HS65_LL_NOR2X6 U14314 ( .A(n2522), .B(n2257), .Z(n2356) );
  HS65_LL_NOR2X6 U14315 ( .A(n1394), .B(n1129), .Z(n1228) );
  HS65_LL_NOR2X6 U14316 ( .A(n1770), .B(n1505), .Z(n1604) );
  HS65_LL_NOR2X6 U14317 ( .A(n2837), .B(n3807), .Z(n3803) );
  HS65_LL_IVX9 U14318 ( .A(n2969), .Z(n631) );
  HS65_LL_NAND2X7 U14319 ( .A(n1180), .B(n1179), .Z(n1185) );
  HS65_LL_IVX9 U14320 ( .A(n1522), .Z(n813) );
  HS65_LL_NOR2X6 U14321 ( .A(n1544), .B(n1537), .Z(n1688) );
  HS65_LL_NOR2X6 U14322 ( .A(n7846), .B(n8106), .Z(n7989) );
  HS65_LL_NOR2X6 U14323 ( .A(n3203), .B(n3197), .Z(n3840) );
  HS65_LL_NOR2X6 U14324 ( .A(n2938), .B(n2931), .Z(n3485) );
  HS65_LL_NOR2X6 U14325 ( .A(n2296), .B(n2289), .Z(n2440) );
  HS65_LL_NOR2X6 U14326 ( .A(n1168), .B(n1161), .Z(n1312) );
  HS65_LL_NOR2X6 U14327 ( .A(n1920), .B(n1913), .Z(n2064) );
  HS65_LL_NOR2X6 U14328 ( .A(n2837), .B(n3183), .Z(n3866) );
  HS65_LL_OAI21X3 U14329 ( .A(n8339), .B(n8369), .C(n8601), .Z(n8890) );
  HS65_LL_NAND4ABX3 U14330 ( .A(n4687), .B(n4688), .C(n4689), .D(n4690), .Z(
        n4544) );
  HS65_LL_NOR4ABX2 U14331 ( .A(n4691), .B(n4692), .C(n4693), .D(n4694), .Z(
        n4690) );
  HS65_LL_NAND4ABX3 U14332 ( .A(n4718), .B(n4719), .C(n4720), .D(n4721), .Z(
        n4688) );
  HS65_LL_MX41X7 U14333 ( .D0(n4481), .S0(n36), .D1(n10), .S1(n42), .D2(n44), 
        .S2(n19), .D3(n39), .S3(n23), .Z(n4687) );
  HS65_LL_NAND4ABX3 U14334 ( .A(n6280), .B(n6281), .C(n6282), .D(n6283), .Z(
        n6137) );
  HS65_LL_NOR4ABX2 U14335 ( .A(n6284), .B(n6285), .C(n6286), .D(n6287), .Z(
        n6283) );
  HS65_LL_NAND4ABX3 U14336 ( .A(n6311), .B(n6312), .C(n6313), .D(n6314), .Z(
        n6281) );
  HS65_LL_MX41X7 U14337 ( .D0(n6074), .S0(n558), .D1(n532), .S1(n564), .D2(
        n566), .S2(n541), .D3(n561), .S3(n545), .Z(n6280) );
  HS65_LL_IVX9 U14338 ( .A(n8238), .Z(n366) );
  HS65_LL_NOR2X6 U14339 ( .A(n1117), .B(n1179), .Z(n1339) );
  HS65_LL_NOR2X6 U14340 ( .A(n1869), .B(n1931), .Z(n2091) );
  HS65_LL_NOR2X6 U14341 ( .A(n2238), .B(n2297), .Z(n2501) );
  HS65_LL_IVX9 U14342 ( .A(n2970), .Z(n651) );
  HS65_LL_NAND4ABX3 U14343 ( .A(n4900), .B(n4901), .C(n4902), .D(n4903), .Z(
        n4742) );
  HS65_LL_NAND4ABX3 U14344 ( .A(n4929), .B(n4930), .C(n4931), .D(n4932), .Z(
        n4901) );
  HS65_LL_NOR4ABX2 U14345 ( .A(n4904), .B(n4905), .C(n4906), .D(n4907), .Z(
        n4903) );
  HS65_LL_MX41X7 U14346 ( .D0(n4589), .S0(n262), .D1(n247), .S1(n264), .D2(
        n255), .S2(n236), .D3(n233), .S3(n268), .Z(n4900) );
  HS65_LL_NAND4ABX3 U14347 ( .A(n4953), .B(n4954), .C(n4955), .D(n4956), .Z(
        n4768) );
  HS65_LL_NAND4ABX3 U14348 ( .A(n4982), .B(n4983), .C(n4984), .D(n4985), .Z(
        n4954) );
  HS65_LL_NOR4ABX2 U14349 ( .A(n4957), .B(n4958), .C(n4959), .D(n4960), .Z(
        n4956) );
  HS65_LL_MX41X7 U14350 ( .D0(n4606), .S0(n479), .D1(n464), .S1(n481), .D2(
        n472), .S2(n453), .D3(n450), .S3(n485), .Z(n4953) );
  HS65_LL_NAND4ABX3 U14351 ( .A(n6546), .B(n6547), .C(n6548), .D(n6549), .Z(
        n6361) );
  HS65_LL_NAND4ABX3 U14352 ( .A(n6575), .B(n6576), .C(n6577), .D(n6578), .Z(
        n6547) );
  HS65_LL_NOR4ABX2 U14353 ( .A(n6550), .B(n6551), .C(n6552), .D(n6553), .Z(
        n6549) );
  HS65_LL_MX41X7 U14354 ( .D0(n6199), .S0(n304), .D1(n289), .S1(n306), .D2(
        n297), .S2(n278), .D3(n275), .S3(n310), .Z(n6546) );
  HS65_LL_NAND4ABX3 U14355 ( .A(n6493), .B(n6494), .C(n6495), .D(n6496), .Z(
        n6322) );
  HS65_LL_NAND4ABX3 U14356 ( .A(n6522), .B(n6523), .C(n6524), .D(n6525), .Z(
        n6494) );
  HS65_LL_NOR4ABX2 U14357 ( .A(n6497), .B(n6498), .C(n6499), .D(n6500), .Z(
        n6496) );
  HS65_LL_MX41X7 U14358 ( .D0(n6182), .S0(n84), .D1(n68), .S1(n78), .D2(n90), 
        .S2(n59), .D3(n64), .S3(n82), .Z(n6493) );
  HS65_LL_NOR2X6 U14359 ( .A(n1862), .B(n1921), .Z(n2125) );
  HS65_LL_NOR2X6 U14360 ( .A(n1110), .B(n1169), .Z(n1373) );
  HS65_LL_NOR2X6 U14361 ( .A(n4448), .B(n4748), .Z(n4929) );
  HS65_LL_NOR2X6 U14362 ( .A(n4509), .B(n4774), .Z(n4982) );
  HS65_LL_NOR2X6 U14363 ( .A(n6102), .B(n6367), .Z(n6575) );
  HS65_LL_NOR2X6 U14364 ( .A(n6041), .B(n6328), .Z(n6522) );
  HS65_LL_NOR2X6 U14365 ( .A(n2245), .B(n2307), .Z(n2467) );
  HS65_LL_IVX9 U14366 ( .A(n7713), .Z(n102) );
  HS65_LL_IVX9 U14367 ( .A(n7675), .Z(n582) );
  HS65_LL_IVX9 U14368 ( .A(n2995), .Z(n442) );
  HS65_LL_IVX9 U14369 ( .A(n2857), .Z(n219) );
  HS65_LL_NOR2X6 U14370 ( .A(n1486), .B(n1545), .Z(n1749) );
  HS65_LL_IVX9 U14371 ( .A(n7767), .Z(n319) );
  HS65_LL_IVX9 U14372 ( .A(n7656), .Z(n122) );
  HS65_LL_IVX9 U14373 ( .A(n7619), .Z(n602) );
  HS65_LL_IVX9 U14374 ( .A(n2257), .Z(n903) );
  HS65_LL_IVX9 U14375 ( .A(n1505), .Z(n821) );
  HS65_LL_IVX9 U14376 ( .A(n1129), .Z(n862) );
  HS65_LL_IVX9 U14377 ( .A(n1881), .Z(n780) );
  HS65_LL_NOR2X6 U14378 ( .A(n1493), .B(n1555), .Z(n1715) );
  HS65_LL_OAI21X3 U14379 ( .A(n2845), .B(n2838), .C(n3355), .Z(n3354) );
  HS65_LL_CBI4I1X5 U14380 ( .A(n7943), .B(n7951), .C(n8363), .D(n8335), .Z(
        n8884) );
  HS65_LL_NOR2X6 U14381 ( .A(n6088), .B(n6569), .Z(n6539) );
  HS65_LL_NOR2X6 U14382 ( .A(n6049), .B(n6516), .Z(n6486) );
  HS65_LL_NOR2X6 U14383 ( .A(n4456), .B(n4923), .Z(n4893) );
  HS65_LL_NOR2X6 U14384 ( .A(n4495), .B(n4976), .Z(n4946) );
  HS65_LL_OAI21X3 U14385 ( .A(n7749), .B(n8082), .C(n8636), .Z(n8635) );
  HS65_LL_CBI4I1X5 U14386 ( .A(n7861), .B(n7850), .C(n8117), .D(n8102), .Z(
        n8944) );
  HS65_LL_IVX9 U14387 ( .A(n5532), .Z(n252) );
  HS65_LL_IVX9 U14388 ( .A(n5554), .Z(n469) );
  HS65_LL_IVX9 U14389 ( .A(n7124), .Z(n89) );
  HS65_LL_IVX9 U14390 ( .A(n7146), .Z(n294) );
  HS65_LL_IVX9 U14391 ( .A(n7171), .Z(n526) );
  HS65_LL_IVX9 U14392 ( .A(n5579), .Z(n702) );
  HS65_LL_NOR2X6 U14393 ( .A(n2889), .B(n3692), .Z(n3688) );
  HS65_LL_NOR2X6 U14394 ( .A(n3972), .B(n2845), .Z(n3375) );
  HS65_LL_NOR2X6 U14395 ( .A(n3952), .B(n2875), .Z(n3321) );
  HS65_LL_NOR2X6 U14396 ( .A(n2069), .B(n1957), .Z(n2124) );
  HS65_LL_NOR2X6 U14397 ( .A(n1317), .B(n1205), .Z(n1372) );
  HS65_LL_CBI4I1X5 U14398 ( .A(n4494), .B(n4603), .C(n4988), .D(n4968), .Z(
        n5903) );
  HS65_LL_CBI4I1X5 U14399 ( .A(n6087), .B(n6196), .C(n6581), .D(n6561), .Z(
        n7495) );
  HS65_LL_CBI4I1X5 U14400 ( .A(n4455), .B(n4586), .C(n4876), .D(n4915), .Z(
        n5844) );
  HS65_LL_CBI4I1X5 U14401 ( .A(n6048), .B(n6179), .C(n6469), .D(n6508), .Z(
        n7436) );
  HS65_LL_IVX9 U14402 ( .A(n2845), .Z(n421) );
  HS65_LL_IVX9 U14403 ( .A(n2875), .Z(n639) );
  HS65_LL_NOR2X6 U14404 ( .A(n1494), .B(n1520), .Z(n1610) );
  HS65_LL_NOR2X6 U14405 ( .A(n2246), .B(n2272), .Z(n2362) );
  HS65_LL_NOR2X6 U14406 ( .A(n1870), .B(n1896), .Z(n1986) );
  HS65_LL_NOR2X6 U14407 ( .A(n1118), .B(n1144), .Z(n1234) );
  HS65_LL_NOR2X6 U14408 ( .A(n2445), .B(n2333), .Z(n2500) );
  HS65_LL_IVX9 U14409 ( .A(n3731), .Z(n625) );
  HS65_LL_IVX9 U14410 ( .A(n7859), .Z(n369) );
  HS65_LL_NOR2X6 U14411 ( .A(n1693), .B(n1581), .Z(n1748) );
  HS65_LL_NOR3X4 U14412 ( .A(n4296), .B(n2849), .C(n3960), .Z(n4293) );
  HS65_LL_OAI21X3 U14413 ( .A(n3197), .B(n3185), .C(n3966), .Z(n4296) );
  HS65_LL_NOR3X4 U14414 ( .A(n4237), .B(n2879), .C(n3940), .Z(n4234) );
  HS65_LL_OAI21X3 U14415 ( .A(n3133), .B(n3158), .C(n3946), .Z(n4237) );
  HS65_LL_IVX9 U14416 ( .A(n3846), .Z(n406) );
  HS65_LL_NAND2X7 U14417 ( .A(n599), .B(n7699), .Z(n8700) );
  HS65_LL_NOR2X6 U14418 ( .A(n4733), .B(n4447), .Z(n5295) );
  HS65_LL_NOR2X6 U14419 ( .A(n6329), .B(n6040), .Z(n6887) );
  HS65_LL_NAND2X7 U14420 ( .A(n612), .B(n7699), .Z(n7791) );
  HS65_LL_NOR2X6 U14421 ( .A(n1931), .B(n1868), .Z(n2040) );
  HS65_LL_NOR2X6 U14422 ( .A(n1179), .B(n1116), .Z(n1288) );
  HS65_LL_IVX9 U14423 ( .A(n1199), .Z(n839) );
  HS65_LL_IVX9 U14424 ( .A(n1951), .Z(n757) );
  HS65_LL_NOR2X6 U14425 ( .A(n2888), .B(n3343), .Z(n3700) );
  HS65_LL_IVX9 U14426 ( .A(n7848), .Z(n396) );
  HS65_LL_IVX9 U14427 ( .A(n4448), .Z(n246) );
  HS65_LL_IVX9 U14428 ( .A(n4509), .Z(n463) );
  HS65_LL_IVX9 U14429 ( .A(n6102), .Z(n288) );
  HS65_LL_IVX9 U14430 ( .A(n6041), .Z(n67) );
  HS65_LL_NOR2X6 U14431 ( .A(n6196), .B(n7221), .Z(n6584) );
  HS65_LL_NOR2X6 U14432 ( .A(n6179), .B(n7196), .Z(n6472) );
  HS65_LL_NOR2X6 U14433 ( .A(n4586), .B(n5604), .Z(n4879) );
  HS65_LL_NOR2X6 U14434 ( .A(n4603), .B(n5629), .Z(n4991) );
  HS65_LL_NOR2X6 U14435 ( .A(n6126), .B(n7170), .Z(n6458) );
  HS65_LL_NOR2X6 U14436 ( .A(n4533), .B(n5578), .Z(n4865) );
  HS65_LL_IVX9 U14437 ( .A(n1493), .Z(n822) );
  HS65_LL_IVX9 U14438 ( .A(n2245), .Z(n904) );
  HS65_LL_IVX9 U14439 ( .A(n1117), .Z(n863) );
  HS65_LL_IVX9 U14440 ( .A(n1869), .Z(n781) );
  HS65_LL_NOR2X6 U14441 ( .A(n3928), .B(n2940), .Z(n3090) );
  HS65_LL_IVX9 U14442 ( .A(n2327), .Z(n880) );
  HS65_LL_NOR2X6 U14443 ( .A(n1555), .B(n1492), .Z(n1664) );
  HS65_LL_NOR2X6 U14444 ( .A(n2307), .B(n2244), .Z(n2416) );
  HS65_LL_NAND2X7 U14445 ( .A(n90), .B(n6182), .Z(n6877) );
  HS65_LL_OAI21X3 U14446 ( .A(n2845), .B(n2846), .C(n2847), .Z(n2844) );
  HS65_LL_OAI21X3 U14447 ( .A(n2940), .B(n3112), .C(n4057), .Z(n4168) );
  HS65_LL_IVX9 U14448 ( .A(n7750), .Z(n367) );
  HS65_LL_IVX9 U14449 ( .A(n1695), .Z(n833) );
  HS65_LL_IVX9 U14450 ( .A(n2447), .Z(n915) );
  HS65_LL_IVX9 U14451 ( .A(n1319), .Z(n874) );
  HS65_LL_IVX9 U14452 ( .A(n2071), .Z(n792) );
  HS65_LL_IVX9 U14453 ( .A(n1575), .Z(n798) );
  HS65_LL_NOR2X6 U14454 ( .A(n2957), .B(n3475), .Z(n3457) );
  HS65_LL_IVX9 U14455 ( .A(n1931), .Z(n770) );
  HS65_LL_IVX9 U14456 ( .A(n1179), .Z(n852) );
  HS65_LL_IVX9 U14457 ( .A(n8117), .Z(n384) );
  HS65_LL_IVX9 U14458 ( .A(n8363), .Z(n345) );
  HS65_LL_IVX9 U14459 ( .A(n4460), .Z(n245) );
  HS65_LL_IVX9 U14460 ( .A(n4499), .Z(n462) );
  HS65_LL_IVX9 U14461 ( .A(n6053), .Z(n69) );
  HS65_LL_IVX9 U14462 ( .A(n6092), .Z(n287) );
  HS65_LL_CBI4I1X5 U14463 ( .A(n8117), .B(n7981), .C(n8238), .D(n8239), .Z(
        n8237) );
  HS65_LL_IVX9 U14464 ( .A(n2119), .Z(n760) );
  HS65_LL_IVX9 U14465 ( .A(n2307), .Z(n893) );
  HS65_LL_OAI21X3 U14466 ( .A(n2875), .B(n2876), .C(n2877), .Z(n2874) );
  HS65_LL_NOR2X6 U14467 ( .A(n7686), .B(n7631), .Z(n8133) );
  HS65_LL_NOR2X6 U14468 ( .A(n7724), .B(n7651), .Z(n8184) );
  HS65_LL_NOR4ABX2 U14469 ( .A(n5899), .B(n5900), .C(n5901), .D(n5902), .Z(
        n5617) );
  HS65_LL_MX41X7 U14470 ( .D0(n454), .S0(n481), .D1(n451), .S1(n485), .D2(n475), .S2(n461), .D3(n478), .S3(n4606), .Z(n5902) );
  HS65_LL_AO212X4 U14471 ( .A(n474), .B(n5430), .C(n473), .D(n452), .E(n5903), 
        .Z(n5901) );
  HS65_LL_NOR3AX2 U14472 ( .A(n5904), .B(n5416), .C(n5460), .Z(n5900) );
  HS65_LL_NOR4ABX2 U14473 ( .A(n7491), .B(n7492), .C(n7493), .D(n7494), .Z(
        n7209) );
  HS65_LL_MX41X7 U14474 ( .D0(n279), .S0(n306), .D1(n276), .S1(n310), .D2(n300), .S2(n286), .D3(n303), .S3(n6199), .Z(n7494) );
  HS65_LL_AO212X4 U14475 ( .A(n299), .B(n7022), .C(n298), .D(n277), .E(n7495), 
        .Z(n7493) );
  HS65_LL_NOR3AX2 U14476 ( .A(n7496), .B(n7008), .C(n7052), .Z(n7492) );
  HS65_LL_NOR4ABX2 U14477 ( .A(n5840), .B(n5841), .C(n5842), .D(n5843), .Z(
        n5592) );
  HS65_LL_MX41X7 U14478 ( .D0(n237), .S0(n264), .D1(n234), .S1(n268), .D2(n258), .S2(n244), .D3(n261), .S3(n4589), .Z(n5843) );
  HS65_LL_AO212X4 U14479 ( .A(n257), .B(n5315), .C(n256), .D(n235), .E(n5844), 
        .Z(n5842) );
  HS65_LL_NOR3AX2 U14480 ( .A(n5845), .B(n5301), .C(n5345), .Z(n5841) );
  HS65_LL_NOR4ABX2 U14481 ( .A(n7432), .B(n7433), .C(n7434), .D(n7435), .Z(
        n7184) );
  HS65_LL_MX41X7 U14482 ( .D0(n58), .S0(n78), .D1(n63), .S1(n82), .D2(n73), 
        .S2(n55), .D3(n85), .S3(n6182), .Z(n7435) );
  HS65_LL_AO212X4 U14483 ( .A(n76), .B(n6907), .C(n74), .D(n66), .E(n7436), 
        .Z(n7434) );
  HS65_LL_NOR3AX2 U14484 ( .A(n7437), .B(n6893), .C(n6937), .Z(n7433) );
  HS65_LL_NOR4ABX2 U14485 ( .A(n5681), .B(n5682), .C(n5683), .D(n5684), .Z(
        n5573) );
  HS65_LL_MX41X7 U14486 ( .D0(n673), .S0(n697), .D1(n679), .S1(n694), .D2(n684), .S2(n670), .D3(n692), .S3(n4521), .Z(n5684) );
  HS65_LL_AO212X4 U14487 ( .A(n688), .B(n5199), .C(n686), .D(n680), .E(n5685), 
        .Z(n5683) );
  HS65_LL_NOR3AX2 U14488 ( .A(n5686), .B(n5185), .C(n5230), .Z(n5682) );
  HS65_LL_NOR4ABX2 U14489 ( .A(n7273), .B(n7274), .C(n7275), .D(n7276), .Z(
        n7165) );
  HS65_LL_MX41X7 U14490 ( .D0(n497), .S0(n521), .D1(n503), .S1(n518), .D2(n508), .S2(n494), .D3(n516), .S3(n6114), .Z(n7276) );
  HS65_LL_AO212X4 U14491 ( .A(n512), .B(n6791), .C(n510), .D(n504), .E(n7277), 
        .Z(n7275) );
  HS65_LL_NOR3AX2 U14492 ( .A(n7278), .B(n6777), .C(n6822), .Z(n7274) );
  HS65_LL_NOR4ABX2 U14493 ( .A(n7243), .B(n7244), .C(n7245), .D(n7246), .Z(
        n7101) );
  HS65_LL_MX41X7 U14494 ( .D0(n540), .S0(n564), .D1(n561), .S1(n546), .D2(n537), .S2(n551), .D3(n559), .S3(n6074), .Z(n7246) );
  HS65_LL_AO212X4 U14495 ( .A(n555), .B(n6670), .C(n553), .D(n547), .E(n7247), 
        .Z(n7245) );
  HS65_LL_NOR3AX2 U14496 ( .A(n7248), .B(n6656), .C(n6687), .Z(n7244) );
  HS65_LL_NOR4ABX2 U14497 ( .A(n5651), .B(n5652), .C(n5653), .D(n5654), .Z(
        n5509) );
  HS65_LL_MX41X7 U14498 ( .D0(n18), .S0(n42), .D1(n39), .S1(n24), .D2(n15), 
        .S2(n29), .D3(n37), .S3(n4481), .Z(n5654) );
  HS65_LL_AO212X4 U14499 ( .A(n33), .B(n5077), .C(n31), .D(n25), .E(n5655), 
        .Z(n5653) );
  HS65_LL_NOR3AX2 U14500 ( .A(n5656), .B(n5063), .C(n5094), .Z(n5652) );
  HS65_LL_NOR3X4 U14501 ( .A(n1433), .B(n1124), .C(n1379), .Z(n1430) );
  HS65_LL_OAI21X3 U14502 ( .A(n1161), .B(n1180), .C(n1388), .Z(n1433) );
  HS65_LL_NOR3X4 U14503 ( .A(n2185), .B(n1876), .C(n2131), .Z(n2182) );
  HS65_LL_OAI21X3 U14504 ( .A(n1913), .B(n1932), .C(n2140), .Z(n2185) );
  HS65_LL_NOR3X4 U14505 ( .A(n1809), .B(n1500), .C(n1755), .Z(n1806) );
  HS65_LL_OAI21X3 U14506 ( .A(n1537), .B(n1556), .C(n1764), .Z(n1809) );
  HS65_LL_NOR3X4 U14507 ( .A(n2561), .B(n2252), .C(n2507), .Z(n2558) );
  HS65_LL_OAI21X3 U14508 ( .A(n2289), .B(n2308), .C(n2516), .Z(n2561) );
  HS65_LL_IVX9 U14509 ( .A(n7831), .Z(n604) );
  HS65_LL_IVX9 U14510 ( .A(n8510), .Z(n323) );
  HS65_LL_IVX9 U14511 ( .A(n4495), .Z(n480) );
  HS65_LL_IVX9 U14512 ( .A(n6088), .Z(n305) );
  HS65_LL_IVX9 U14513 ( .A(n4456), .Z(n263) );
  HS65_LL_IVX9 U14514 ( .A(n6049), .Z(n86) );
  HS65_LL_IVX9 U14515 ( .A(n6588), .Z(n301) );
  HS65_LL_IVX9 U14516 ( .A(n6476), .Z(n77) );
  HS65_LL_IVX9 U14517 ( .A(n4995), .Z(n476) );
  HS65_LL_IVX9 U14518 ( .A(n1555), .Z(n811) );
  HS65_LL_IVX9 U14519 ( .A(n5507), .Z(n35) );
  HS65_LL_IVX9 U14520 ( .A(n7099), .Z(n557) );
  HS65_LL_IVX9 U14521 ( .A(n2495), .Z(n883) );
  HS65_LL_IVX9 U14522 ( .A(n1367), .Z(n842) );
  HS65_LL_IVX9 U14523 ( .A(n1743), .Z(n801) );
  HS65_LL_NOR2X6 U14524 ( .A(n2307), .B(n2273), .Z(n2499) );
  HS65_LL_NOR2X6 U14525 ( .A(n1555), .B(n1521), .Z(n1747) );
  HS65_LL_NOR2X6 U14526 ( .A(n1931), .B(n1897), .Z(n2123) );
  HS65_LL_NOR2X6 U14527 ( .A(n1179), .B(n1145), .Z(n1371) );
  HS65_LL_IVX9 U14528 ( .A(n5533), .Z(n260) );
  HS65_LL_IVX9 U14529 ( .A(n5555), .Z(n477) );
  HS65_LL_IVX9 U14530 ( .A(n5571), .Z(n690) );
  HS65_LL_IVX9 U14531 ( .A(n7125), .Z(n83) );
  HS65_LL_IVX9 U14532 ( .A(n7147), .Z(n302) );
  HS65_LL_IVX9 U14533 ( .A(n7163), .Z(n514) );
  HS65_LL_NOR2X6 U14534 ( .A(n7846), .B(n7860), .Z(n8276) );
  HS65_LL_IVX9 U14535 ( .A(n8556), .Z(n326) );
  HS65_LL_NAND2X7 U14536 ( .A(n2447), .B(n2273), .Z(n2388) );
  HS65_LL_NAND2X7 U14537 ( .A(n1695), .B(n1521), .Z(n1636) );
  HS65_LL_NOR4ABX2 U14538 ( .A(n3336), .B(n3337), .C(n3338), .D(n3339), .Z(
        n2975) );
  HS65_LL_OAI222X2 U14539 ( .A(n3342), .B(n3343), .C(n2889), .D(n2881), .E(
        n3133), .F(n3129), .Z(n3338) );
  HS65_LL_NOR3X4 U14540 ( .A(n3344), .B(n3345), .C(n3346), .Z(n3337) );
  HS65_LL_OAI212X5 U14541 ( .A(n3340), .B(n2876), .C(n3128), .D(n2890), .E(
        n3341), .Z(n3339) );
  HS65_LL_NAND2X7 U14542 ( .A(n1319), .B(n1145), .Z(n1260) );
  HS65_LL_NAND2X7 U14543 ( .A(n2071), .B(n1897), .Z(n2012) );
  HS65_LL_IVX9 U14544 ( .A(n3491), .Z(n203) );
  HS65_LL_OAI21X3 U14545 ( .A(n7767), .B(n8357), .C(n8621), .Z(n8620) );
  HS65_LL_NAND2X7 U14546 ( .A(n3846), .B(n2994), .Z(n3775) );
  HS65_LL_IVX9 U14547 ( .A(n8106), .Z(n398) );
  HS65_LL_NOR2X6 U14548 ( .A(n7980), .B(n7847), .Z(n8305) );
  HS65_LL_NOR2X6 U14549 ( .A(n7850), .B(n8649), .Z(n8120) );
  HS65_LL_NAND2X7 U14550 ( .A(n8254), .B(n7847), .Z(n8195) );
  HS65_LL_IVX9 U14551 ( .A(n1863), .Z(n759) );
  HS65_LL_NOR4ABX2 U14552 ( .A(n5543), .B(n5551), .C(n4513), .D(n5615), .Z(
        n5614) );
  HS65_LL_OAI212X5 U14553 ( .A(n5555), .B(n4494), .C(n5616), .D(n4499), .E(
        n5617), .Z(n5615) );
  HS65_LL_NOR4ABX2 U14554 ( .A(n7135), .B(n7143), .C(n6106), .D(n7207), .Z(
        n7206) );
  HS65_LL_OAI212X5 U14555 ( .A(n7147), .B(n6087), .C(n7208), .D(n6092), .E(
        n7209), .Z(n7207) );
  HS65_LL_NOR4ABX2 U14556 ( .A(n7079), .B(n7160), .C(n7161), .D(n7162), .Z(
        n7159) );
  HS65_LL_OAI212X5 U14557 ( .A(n7163), .B(n6219), .C(n7164), .D(n6118), .E(
        n7165), .Z(n7162) );
  HS65_LL_NOR4ABX2 U14558 ( .A(n5487), .B(n5568), .C(n5569), .D(n5570), .Z(
        n5567) );
  HS65_LL_OAI212X5 U14559 ( .A(n5571), .B(n4626), .C(n5572), .D(n4525), .E(
        n5573), .Z(n5570) );
  HS65_LL_CBI4I1X5 U14560 ( .A(n1317), .B(n1109), .C(n1161), .D(n1420), .Z(
        n1398) );
  HS65_LL_AO12X9 U14561 ( .A(n1168), .B(n1149), .C(n1369), .Z(n1420) );
  HS65_LL_CBI4I1X5 U14562 ( .A(n2069), .B(n1861), .C(n1913), .D(n2172), .Z(
        n2150) );
  HS65_LL_AO12X9 U14563 ( .A(n1920), .B(n1901), .C(n2121), .Z(n2172) );
  HS65_LL_IVX9 U14564 ( .A(n4747), .Z(n261) );
  HS65_LL_IVX9 U14565 ( .A(n4773), .Z(n478) );
  HS65_LL_IVX9 U14566 ( .A(n6327), .Z(n85) );
  HS65_LL_IVX9 U14567 ( .A(n6366), .Z(n303) );
  HS65_LL_CBI4I1X5 U14568 ( .A(n2445), .B(n2237), .C(n2289), .D(n2548), .Z(
        n2526) );
  HS65_LL_AO12X9 U14569 ( .A(n2296), .B(n2277), .C(n2497), .Z(n2548) );
  HS65_LL_NOR2X6 U14570 ( .A(n2273), .B(n2520), .Z(n2293) );
  HS65_LL_IVX9 U14571 ( .A(n7941), .Z(n332) );
  HS65_LL_IVX9 U14572 ( .A(n7835), .Z(n578) );
  HS65_LL_IVX9 U14573 ( .A(n7874), .Z(n98) );
  HS65_LL_NOR2X6 U14574 ( .A(n8048), .B(n7948), .Z(n8519) );
  HS65_LL_IVX9 U14575 ( .A(n1111), .Z(n841) );
  HS65_LL_IVX9 U14576 ( .A(n1487), .Z(n800) );
  HS65_LL_IVX9 U14577 ( .A(n2239), .Z(n882) );
  HS65_LL_NOR2X6 U14578 ( .A(n7993), .B(n8238), .Z(n8208) );
  HS65_LL_NOR2X6 U14579 ( .A(n1897), .B(n2144), .Z(n1917) );
  HS65_LL_NOR2X6 U14580 ( .A(n1145), .B(n1392), .Z(n1165) );
  HS65_LL_NOR2X6 U14581 ( .A(n8449), .B(n7663), .Z(n8185) );
  HS65_LL_IVX9 U14582 ( .A(n7980), .Z(n399) );
  HS65_LL_IVX9 U14583 ( .A(n8048), .Z(n350) );
  HS65_LL_IVX9 U14584 ( .A(n7624), .Z(n591) );
  HS65_LL_IVX9 U14585 ( .A(n7664), .Z(n111) );
  HS65_LL_NOR2X6 U14586 ( .A(n1521), .B(n1768), .Z(n1541) );
  HS65_LL_NAND2X7 U14587 ( .A(n3731), .B(n2969), .Z(n3660) );
  HS65_LL_OAI21X3 U14588 ( .A(n1957), .B(n1863), .C(n2021), .Z(n2200) );
  HS65_LL_IVX9 U14589 ( .A(n8058), .Z(n352) );
  HS65_LL_NOR2X6 U14590 ( .A(n2994), .B(n3970), .Z(n3200) );
  HS65_LL_NOR2X6 U14591 ( .A(n2856), .B(n3926), .Z(n2935) );
  HS65_LL_NOR2X6 U14592 ( .A(n6859), .B(n6040), .Z(n6879) );
  HS65_LL_IVX9 U14593 ( .A(n7949), .Z(n356) );
  HS65_LL_NOR4ABX2 U14594 ( .A(n3961), .B(n3962), .C(n3963), .D(n3964), .Z(
        n2848) );
  HS65_LL_CBI4I1X5 U14595 ( .A(n2845), .B(n3412), .C(n2995), .D(n3372), .Z(
        n3963) );
  HS65_LL_CBI4I1X5 U14596 ( .A(n3832), .B(n3204), .C(n2836), .D(n3965), .Z(
        n3964) );
  HS65_LL_NOR4ABX2 U14597 ( .A(n3785), .B(n3837), .C(n3857), .D(n3880), .Z(
        n3961) );
  HS65_LL_OAI21X3 U14598 ( .A(n1205), .B(n1111), .C(n1269), .Z(n1448) );
  HS65_LL_OAI21X3 U14599 ( .A(n1581), .B(n1487), .C(n1645), .Z(n1824) );
  HS65_LL_OAI21X3 U14600 ( .A(n2333), .B(n2239), .C(n2397), .Z(n2576) );
  HS65_LL_NOR4ABX2 U14601 ( .A(n7936), .B(n7937), .C(n7938), .D(n7939), .Z(
        n7935) );
  HS65_LL_OAI212X5 U14602 ( .A(n7940), .B(n7941), .C(n7942), .D(n7943), .E(
        n7944), .Z(n7938) );
  HS65_LL_IVX9 U14603 ( .A(n3342), .Z(n633) );
  HS65_LL_NOR2X6 U14604 ( .A(n3450), .B(n3491), .Z(n3458) );
  HS65_LL_NOR4ABX2 U14605 ( .A(n4186), .B(n4187), .C(n4188), .D(n4189), .Z(
        n3896) );
  HS65_LL_CBI4I1X5 U14606 ( .A(n2940), .B(n3067), .C(n2857), .D(n3087), .Z(
        n4188) );
  HS65_LL_CBI4I1X5 U14607 ( .A(n3477), .B(n2939), .C(n3475), .D(n4190), .Z(
        n4189) );
  HS65_LL_NOR4ABX2 U14608 ( .A(n3427), .B(n3482), .C(n3502), .D(n3526), .Z(
        n4186) );
  HS65_LL_OAI21X3 U14609 ( .A(n2875), .B(n2890), .C(n3301), .Z(n3300) );
  HS65_LL_NOR2X6 U14610 ( .A(n2972), .B(n3950), .Z(n3296) );
  HS65_LL_NOR2X6 U14611 ( .A(n2969), .B(n3950), .Z(n3137) );
  HS65_LL_NOR4ABX2 U14612 ( .A(n3957), .B(n3958), .C(n3959), .D(n3960), .Z(
        n3956) );
  HS65_LL_OAI212X5 U14613 ( .A(n3406), .B(n3396), .C(n3185), .D(n2832), .E(
        n2848), .Z(n3959) );
  HS65_LL_IVX9 U14614 ( .A(n3692), .Z(n661) );
  HS65_LL_NAND4ABX3 U14615 ( .A(n8851), .B(n8852), .C(n8853), .D(n8854), .Z(
        n8622) );
  HS65_LL_NOR4ABX2 U14616 ( .A(n8602), .B(n8588), .C(n8549), .D(n8566), .Z(
        n8853) );
  HS65_LL_CB4I6X9 U14617 ( .A(n319), .B(n329), .C(n356), .D(n8334), .Z(n8851)
         );
  HS65_LL_CBI4I1X5 U14618 ( .A(n8542), .B(n8039), .C(n8540), .D(n8863), .Z(
        n8852) );
  HS65_LL_NAND4ABX3 U14619 ( .A(n8638), .B(n8639), .C(n8640), .D(n8641), .Z(
        n8485) );
  HS65_LL_CB4I6X9 U14620 ( .A(n365), .B(n377), .C(n396), .D(n8101), .Z(n8638)
         );
  HS65_LL_CBI4I1X5 U14621 ( .A(n8240), .B(n7971), .C(n8238), .D(n8651), .Z(
        n8639) );
  HS65_LL_NOR4ABX2 U14622 ( .A(n8221), .B(n8245), .C(n8264), .D(n8287), .Z(
        n8640) );
  HS65_LL_NAND4ABX3 U14623 ( .A(n5546), .B(n5547), .C(n5548), .D(n5549), .Z(
        n4511) );
  HS65_LL_CB4I6X9 U14624 ( .A(n463), .B(n449), .C(n476), .D(n4981), .Z(n5546)
         );
  HS65_LL_NOR4ABX2 U14625 ( .A(n5381), .B(n5399), .C(n5457), .D(n5413), .Z(
        n5548) );
  HS65_LL_CBI4I1X5 U14626 ( .A(n5367), .B(n5555), .C(n4499), .D(n5556), .Z(
        n5547) );
  HS65_LL_NAND4ABX3 U14627 ( .A(n5524), .B(n5525), .C(n5526), .D(n5527), .Z(
        n4450) );
  HS65_LL_CB4I6X9 U14628 ( .A(n246), .B(n232), .C(n259), .D(n4928), .Z(n5524)
         );
  HS65_LL_NOR4ABX2 U14629 ( .A(n5266), .B(n5284), .C(n5342), .D(n5298), .Z(
        n5526) );
  HS65_LL_CBI4I1X5 U14630 ( .A(n5252), .B(n5533), .C(n4460), .D(n5534), .Z(
        n5525) );
  HS65_LL_NAND4ABX3 U14631 ( .A(n7138), .B(n7139), .C(n7140), .D(n7141), .Z(
        n6104) );
  HS65_LL_CB4I6X9 U14632 ( .A(n288), .B(n274), .C(n301), .D(n6574), .Z(n7138)
         );
  HS65_LL_NOR4ABX2 U14633 ( .A(n6973), .B(n6991), .C(n7049), .D(n7005), .Z(
        n7140) );
  HS65_LL_CBI4I1X5 U14634 ( .A(n6959), .B(n7147), .C(n6092), .D(n7148), .Z(
        n7139) );
  HS65_LL_NAND4ABX3 U14635 ( .A(n9058), .B(n9059), .C(n9060), .D(n9061), .Z(
        n7899) );
  HS65_LL_CB4I6X9 U14636 ( .A(n102), .B(n108), .C(n136), .D(n8452), .Z(n9058)
         );
  HS65_LL_CBI4I1X5 U14637 ( .A(n8767), .B(n7651), .C(n7652), .D(n9079), .Z(
        n9059) );
  HS65_LL_NOR4ABX2 U14638 ( .A(n8778), .B(n8789), .C(n8816), .D(n8800), .Z(
        n9060) );
  HS65_LL_NAND4ABX3 U14639 ( .A(n5779), .B(n5780), .C(n5781), .D(n5782), .Z(
        n5490) );
  HS65_LL_CB4I6X9 U14640 ( .A(n668), .B(n677), .C(n685), .D(n4855), .Z(n5779)
         );
  HS65_LL_NOR4ABX2 U14641 ( .A(n5149), .B(n5167), .C(n5227), .D(n5182), .Z(
        n5781) );
  HS65_LL_CBI4I1X5 U14642 ( .A(n5134), .B(n5571), .C(n4525), .D(n5811), .Z(
        n5780) );
  HS65_LL_NAND4ABX3 U14643 ( .A(n9000), .B(n9001), .C(n9002), .D(n9003), .Z(
        n7800) );
  HS65_LL_CB4I6X9 U14644 ( .A(n582), .B(n588), .C(n616), .D(n8400), .Z(n9000)
         );
  HS65_LL_CBI4I1X5 U14645 ( .A(n8677), .B(n7631), .C(n7632), .D(n9021), .Z(
        n9001) );
  HS65_LL_NOR4ABX2 U14646 ( .A(n8688), .B(n8699), .C(n8726), .D(n8710), .Z(
        n9002) );
  HS65_LL_NAND4ABX3 U14647 ( .A(n7371), .B(n7372), .C(n7373), .D(n7374), .Z(
        n7082) );
  HS65_LL_CB4I6X9 U14648 ( .A(n492), .B(n501), .C(n509), .D(n6448), .Z(n7371)
         );
  HS65_LL_NOR4ABX2 U14649 ( .A(n6741), .B(n6759), .C(n6819), .D(n6774), .Z(
        n7373) );
  HS65_LL_CBI4I1X5 U14650 ( .A(n6726), .B(n7163), .C(n6118), .D(n7403), .Z(
        n7372) );
  HS65_LL_NAND4ABX3 U14651 ( .A(n7116), .B(n7117), .C(n7118), .D(n7119), .Z(
        n6043) );
  HS65_LL_CB4I6X9 U14652 ( .A(n67), .B(n65), .C(n77), .D(n6521), .Z(n7116) );
  HS65_LL_NOR4ABX2 U14653 ( .A(n6858), .B(n6876), .C(n6934), .D(n6890), .Z(
        n7118) );
  HS65_LL_CBI4I1X5 U14654 ( .A(n6844), .B(n7125), .C(n6053), .D(n7126), .Z(
        n7117) );
  HS65_LL_NAND4ABX3 U14655 ( .A(n5717), .B(n5718), .C(n5719), .D(n5720), .Z(
        n5476) );
  HS65_LL_CB4I6X9 U14656 ( .A(n11), .B(n22), .C(n30), .D(n4717), .Z(n5717) );
  HS65_LL_NOR4ABX2 U14657 ( .A(n5027), .B(n5045), .C(n5091), .D(n5060), .Z(
        n5719) );
  HS65_LL_CBI4I1X5 U14658 ( .A(n5012), .B(n5507), .C(n4485), .D(n5749), .Z(
        n5718) );
  HS65_LL_NAND4ABX3 U14659 ( .A(n7309), .B(n7310), .C(n7311), .D(n7312), .Z(
        n7068) );
  HS65_LL_CB4I6X9 U14660 ( .A(n533), .B(n544), .C(n552), .D(n6310), .Z(n7309)
         );
  HS65_LL_NOR4ABX2 U14661 ( .A(n6620), .B(n6638), .C(n6684), .D(n6653), .Z(
        n7311) );
  HS65_LL_CBI4I1X5 U14662 ( .A(n6605), .B(n7099), .C(n6078), .D(n7341), .Z(
        n7310) );
  HS65_LL_CBI4I1X5 U14663 ( .A(n1144), .B(n1145), .C(n1146), .D(n1147), .Z(
        n1134) );
  HS65_LL_OAI21X3 U14664 ( .A(n840), .B(n855), .C(n868), .Z(n1147) );
  HS65_LL_OAI21X3 U14665 ( .A(n3412), .B(n2831), .C(n3784), .Z(n4311) );
  HS65_LL_IVX9 U14666 ( .A(n7861), .Z(n363) );
  HS65_LL_NOR4ABX2 U14667 ( .A(n3941), .B(n3942), .C(n3943), .D(n3944), .Z(
        n2878) );
  HS65_LL_CBI4I1X5 U14668 ( .A(n2875), .B(n3299), .C(n2970), .D(n3318), .Z(
        n3943) );
  HS65_LL_CBI4I1X5 U14669 ( .A(n3717), .B(n3141), .C(n2888), .D(n3945), .Z(
        n3944) );
  HS65_LL_NOR4ABX2 U14670 ( .A(n3670), .B(n3723), .C(n3742), .D(n3765), .Z(
        n3941) );
  HS65_LL_NOR2X6 U14671 ( .A(n8369), .B(n8058), .Z(n8520) );
  HS65_LL_IVX9 U14672 ( .A(n8254), .Z(n372) );
  HS65_LL_IVX9 U14673 ( .A(n3140), .Z(n645) );
  HS65_LL_IVX9 U14674 ( .A(n8123), .Z(n377) );
  HS65_LL_IVX9 U14675 ( .A(n8369), .Z(n329) );
  HS65_LL_OAI21X3 U14676 ( .A(n3299), .B(n2883), .C(n3669), .Z(n4252) );
  HS65_LL_NOR2X6 U14677 ( .A(n1233), .B(n1168), .Z(n1182) );
  HS65_LL_IVX9 U14678 ( .A(n7768), .Z(n333) );
  HS65_LL_NOR4ABX2 U14679 ( .A(n3957), .B(n4024), .C(n2850), .D(n4025), .Z(
        n4023) );
  HS65_LL_OA212X4 U14680 ( .A(n2832), .B(n3204), .C(n3807), .D(n2836), .E(
        n3967), .Z(n4024) );
  HS65_LL_IVX9 U14681 ( .A(n2997), .Z(n408) );
  HS65_LL_IVX9 U14682 ( .A(n2972), .Z(n627) );
  HS65_LL_IVX9 U14683 ( .A(n2859), .Z(n202) );
  HS65_LL_OAI21X3 U14684 ( .A(n3067), .B(n3095), .C(n3426), .Z(n4208) );
  HS65_LL_NOR4ABX2 U14685 ( .A(n7646), .B(n7647), .C(n7648), .D(n7649), .Z(
        n7645) );
  HS65_LL_OA212X4 U14686 ( .A(n7650), .B(n7651), .C(n7652), .D(n7653), .E(
        n7654), .Z(n7647) );
  HS65_LL_OAI21X3 U14687 ( .A(n8106), .B(n8123), .C(n8220), .Z(n8950) );
  HS65_LL_IVX9 U14688 ( .A(n3116), .Z(n193) );
  HS65_LL_IVX9 U14689 ( .A(n2837), .Z(n418) );
  HS65_LL_IVX9 U14690 ( .A(n2889), .Z(n636) );
  HS65_LL_IVX9 U14691 ( .A(n7942), .Z(n344) );
  HS65_LL_IVX9 U14692 ( .A(n3807), .Z(n430) );
  HS65_LL_OAI212X5 U14693 ( .A(n8905), .B(n8540), .C(n8058), .D(n8510), .E(
        n8906), .Z(n8904) );
  HS65_LL_OAI21X3 U14694 ( .A(n330), .B(n334), .C(n341), .Z(n8906) );
  HS65_LL_NOR3X4 U14695 ( .A(n349), .B(n347), .C(n348), .Z(n8905) );
  HS65_LL_IVX9 U14696 ( .A(n7860), .Z(n383) );
  HS65_LL_IVX9 U14697 ( .A(n7769), .Z(n342) );
  HS65_LL_IVX9 U14698 ( .A(n3203), .Z(n432) );
  HS65_LL_IVX9 U14699 ( .A(n2832), .Z(n422) );
  HS65_LL_NOR3AX2 U14700 ( .A(n4057), .B(n4058), .C(n3894), .Z(n4054) );
  HS65_LL_OAI21X3 U14701 ( .A(n2931), .B(n2958), .C(n4064), .Z(n4058) );
  HS65_LL_IVX9 U14702 ( .A(n3299), .Z(n628) );
  HS65_LL_IVX9 U14703 ( .A(n7686), .Z(n590) );
  HS65_LL_NAND2X7 U14704 ( .A(n561), .B(n6074), .Z(n6645) );
  HS65_LL_NAND2X7 U14705 ( .A(n39), .B(n4481), .Z(n5052) );
  HS65_LL_NAND2X7 U14706 ( .A(n600), .B(n7699), .Z(n8392) );
  HS65_LL_IVX9 U14707 ( .A(n8649), .Z(n394) );
  HS65_LL_IVX9 U14708 ( .A(n7971), .Z(n400) );
  HS65_LL_OAI212X5 U14709 ( .A(n4030), .B(n2836), .C(n3397), .D(n2992), .E(
        n4031), .Z(n4029) );
  HS65_LL_OAI21X3 U14710 ( .A(n413), .B(n417), .C(n429), .Z(n4031) );
  HS65_LL_NOR3X4 U14711 ( .A(n439), .B(n435), .C(n431), .Z(n4030) );
  HS65_LL_OAI212X5 U14712 ( .A(n4178), .B(n3475), .C(n3115), .D(n3464), .E(
        n4179), .Z(n4177) );
  HS65_LL_OAI21X3 U14713 ( .A(n198), .B(n194), .C(n210), .Z(n4179) );
  HS65_LL_NOR3X4 U14714 ( .A(n213), .B(n223), .C(n225), .Z(n4178) );
  HS65_LL_IVX9 U14715 ( .A(n4477), .Z(n21) );
  HS65_LL_IVX9 U14716 ( .A(n6070), .Z(n543) );
  HS65_LL_IVX9 U14717 ( .A(n3326), .Z(n630) );
  HS65_LL_IVX9 U14718 ( .A(n4566), .Z(n17) );
  HS65_LL_IVX9 U14719 ( .A(n6159), .Z(n539) );
  HS65_LL_NOR2X6 U14720 ( .A(n8173), .B(n7714), .Z(n8807) );
  HS65_LL_NOR2X6 U14721 ( .A(n8527), .B(n8556), .Z(n8512) );
  HS65_LL_NAND2X7 U14722 ( .A(n518), .B(n6114), .Z(n6766) );
  HS65_LL_NAND2X7 U14723 ( .A(n694), .B(n4521), .Z(n5174) );
  HS65_LL_NAND2X7 U14724 ( .A(n253), .B(n4589), .Z(n4914) );
  HS65_LL_NAND2X7 U14725 ( .A(n470), .B(n4606), .Z(n4967) );
  HS65_LL_NAND2X7 U14726 ( .A(n295), .B(n6199), .Z(n6560) );
  HS65_LL_NAND2X7 U14727 ( .A(n88), .B(n6182), .Z(n6507) );
  HS65_LL_NAND2X7 U14728 ( .A(n485), .B(n4606), .Z(n5405) );
  HS65_LL_NAND2X7 U14729 ( .A(n268), .B(n4589), .Z(n5290) );
  HS65_LL_NAND2X7 U14730 ( .A(n310), .B(n6199), .Z(n6997) );
  HS65_LL_NAND2X7 U14731 ( .A(n82), .B(n6182), .Z(n6882) );
  HS65_LL_IVX9 U14732 ( .A(n4710), .Z(n24) );
  HS65_LL_IVX9 U14733 ( .A(n6303), .Z(n546) );
  HS65_LL_IVX9 U14734 ( .A(n3412), .Z(n409) );
  HS65_LL_IVX9 U14735 ( .A(n7992), .Z(n376) );
  HS65_LL_IVX9 U14736 ( .A(n1168), .Z(n853) );
  HS65_LL_IVX9 U14737 ( .A(n1920), .Z(n771) );
  HS65_LL_IVX9 U14738 ( .A(n2836), .Z(n420) );
  HS65_LL_IVX9 U14739 ( .A(n2273), .Z(n907) );
  HS65_LL_IVX9 U14740 ( .A(n1521), .Z(n825) );
  HS65_LL_IVX9 U14741 ( .A(n1145), .Z(n866) );
  HS65_LL_IVX9 U14742 ( .A(n1897), .Z(n784) );
  HS65_LL_IVX9 U14743 ( .A(n8630), .Z(n354) );
  HS65_LL_IVX9 U14744 ( .A(n2994), .Z(n413) );
  HS65_LL_IVX9 U14745 ( .A(n2296), .Z(n894) );
  HS65_LL_IVX9 U14746 ( .A(n7948), .Z(n330) );
  HS65_LL_NOR2X6 U14747 ( .A(n3140), .B(n3128), .Z(n3662) );
  HS65_LL_OAI21X3 U14748 ( .A(n1367), .B(n1198), .C(n1427), .Z(n1426) );
  HS65_LL_OAI21X3 U14749 ( .A(n862), .B(n865), .C(n847), .Z(n1427) );
  HS65_LL_NAND4ABX3 U14750 ( .A(n4910), .B(n4911), .C(n4912), .D(n4913), .Z(
        n4581) );
  HS65_LL_OAI222X2 U14751 ( .A(n4922), .B(n4456), .C(n4923), .D(n4748), .E(
        n4453), .F(n4448), .Z(n4911) );
  HS65_LL_NOR4ABX2 U14752 ( .A(n4914), .B(n4915), .C(n4916), .D(n4917), .Z(
        n4913) );
  HS65_LL_NAND3X5 U14753 ( .A(n4924), .B(n4925), .C(n4926), .Z(n4910) );
  HS65_LL_NAND4ABX3 U14754 ( .A(n6556), .B(n6557), .C(n6558), .D(n6559), .Z(
        n6191) );
  HS65_LL_OAI222X2 U14755 ( .A(n6568), .B(n6088), .C(n6569), .D(n6367), .E(
        n6085), .F(n6102), .Z(n6557) );
  HS65_LL_NOR4ABX2 U14756 ( .A(n6560), .B(n6561), .C(n6562), .D(n6563), .Z(
        n6559) );
  HS65_LL_NAND3X5 U14757 ( .A(n6570), .B(n6571), .C(n6572), .Z(n6556) );
  HS65_LL_NAND4ABX3 U14758 ( .A(n6503), .B(n6504), .C(n6505), .D(n6506), .Z(
        n6174) );
  HS65_LL_OAI222X2 U14759 ( .A(n6515), .B(n6049), .C(n6516), .D(n6328), .E(
        n6046), .F(n6041), .Z(n6504) );
  HS65_LL_NOR4ABX2 U14760 ( .A(n6507), .B(n6508), .C(n6509), .D(n6510), .Z(
        n6506) );
  HS65_LL_NAND3X5 U14761 ( .A(n6517), .B(n6518), .C(n6519), .Z(n6503) );
  HS65_LL_NOR2X6 U14762 ( .A(n1110), .B(n1168), .Z(n1264) );
  HS65_LL_NOR2X6 U14763 ( .A(n8254), .B(n7860), .Z(n8255) );
  HS65_LL_IVX9 U14764 ( .A(n1544), .Z(n812) );
  HS65_LL_IVX9 U14765 ( .A(n4922), .Z(n234) );
  HS65_LL_IVX9 U14766 ( .A(n6568), .Z(n276) );
  HS65_LL_IVX9 U14767 ( .A(n6515), .Z(n63) );
  HS65_LL_IVX9 U14768 ( .A(n4975), .Z(n451) );
  HS65_LL_NOR2X6 U14769 ( .A(n1199), .B(n1205), .Z(n1120) );
  HS65_LL_OAI21X3 U14770 ( .A(n6094), .B(n6102), .C(n6531), .Z(n6530) );
  HS65_LL_OAI21X3 U14771 ( .A(n6055), .B(n6041), .C(n6478), .Z(n6477) );
  HS65_LL_OAI21X3 U14772 ( .A(n4462), .B(n4448), .C(n4885), .Z(n4884) );
  HS65_LL_IVX9 U14773 ( .A(n3141), .Z(n653) );
  HS65_LL_OAI21X3 U14774 ( .A(n4508), .B(n4509), .C(n4510), .Z(n4507) );
  HS65_LL_OAI21X3 U14775 ( .A(n6101), .B(n6102), .C(n6103), .Z(n6100) );
  HS65_LL_IVX9 U14776 ( .A(n7714), .Z(n129) );
  HS65_LL_IVX9 U14777 ( .A(n7676), .Z(n609) );
  HS65_LL_IVX9 U14778 ( .A(n7943), .Z(n320) );
  HS65_LL_IVX9 U14779 ( .A(n6179), .Z(n62) );
  HS65_LL_IVX9 U14780 ( .A(n4586), .Z(n240) );
  HS65_LL_IVX9 U14781 ( .A(n4603), .Z(n457) );
  HS65_LL_IVX9 U14782 ( .A(n4533), .Z(n676) );
  HS65_LL_IVX9 U14783 ( .A(n6196), .Z(n282) );
  HS65_LL_IVX9 U14784 ( .A(n6126), .Z(n500) );
  HS65_LL_IVX9 U14785 ( .A(n2856), .Z(n198) );
  HS65_LL_NAND4ABX3 U14786 ( .A(n4124), .B(n4125), .C(n4126), .D(n4127), .Z(
        n3910) );
  HS65_LL_CBI4I1X5 U14787 ( .A(n3225), .B(n3286), .C(n2915), .D(n3550), .Z(
        n4124) );
  HS65_LL_NOR4ABX2 U14788 ( .A(n3629), .B(n3653), .C(n3611), .D(n3254), .Z(
        n4126) );
  HS65_LL_CBI4I1X5 U14789 ( .A(n3601), .B(n3994), .C(n3053), .D(n4156), .Z(
        n4125) );
  HS65_LL_NAND4ABX3 U14790 ( .A(n1305), .B(n1306), .C(n1307), .D(n1308), .Z(
        n1174) );
  HS65_LL_NOR3X4 U14791 ( .A(n1313), .B(n1314), .C(n1315), .Z(n1307) );
  HS65_LL_OAI212X5 U14792 ( .A(n1316), .B(n1317), .C(n1146), .D(n1110), .E(
        n1318), .Z(n1306) );
  HS65_LL_NOR4ABX2 U14793 ( .A(n1309), .B(n1310), .C(n1311), .D(n1312), .Z(
        n1308) );
  HS65_LL_NAND4ABX3 U14794 ( .A(n2057), .B(n2058), .C(n2059), .D(n2060), .Z(
        n1926) );
  HS65_LL_NOR3X4 U14795 ( .A(n2065), .B(n2066), .C(n2067), .Z(n2059) );
  HS65_LL_OAI212X5 U14796 ( .A(n2068), .B(n2069), .C(n1898), .D(n1862), .E(
        n2070), .Z(n2058) );
  HS65_LL_NOR4ABX2 U14797 ( .A(n2061), .B(n2062), .C(n2063), .D(n2064), .Z(
        n2060) );
  HS65_LL_NAND4ABX3 U14798 ( .A(n2433), .B(n2434), .C(n2435), .D(n2436), .Z(
        n2302) );
  HS65_LL_NOR3X4 U14799 ( .A(n2441), .B(n2442), .C(n2443), .Z(n2435) );
  HS65_LL_OAI212X5 U14800 ( .A(n2444), .B(n2445), .C(n2274), .D(n2238), .E(
        n2446), .Z(n2434) );
  HS65_LL_NOR4ABX2 U14801 ( .A(n2437), .B(n2438), .C(n2439), .D(n2440), .Z(
        n2436) );
  HS65_LL_NAND4ABX3 U14802 ( .A(n3833), .B(n3834), .C(n3835), .D(n3836), .Z(
        n3169) );
  HS65_LL_NOR3X4 U14803 ( .A(n3841), .B(n3842), .C(n3843), .Z(n3835) );
  HS65_LL_NAND4ABX3 U14804 ( .A(n3847), .B(n3848), .C(n3849), .D(n3850), .Z(
        n3833) );
  HS65_LL_OAI212X5 U14805 ( .A(n3844), .B(n3397), .C(n2995), .D(n2830), .E(
        n3845), .Z(n3834) );
  HS65_LL_NAND4ABX3 U14806 ( .A(n1681), .B(n1682), .C(n1683), .D(n1684), .Z(
        n1550) );
  HS65_LL_NOR3X4 U14807 ( .A(n1689), .B(n1690), .C(n1691), .Z(n1683) );
  HS65_LL_OAI212X5 U14808 ( .A(n1692), .B(n1693), .C(n1522), .D(n1486), .E(
        n1694), .Z(n1682) );
  HS65_LL_NAND4ABX3 U14809 ( .A(n1696), .B(n1697), .C(n1698), .D(n1699), .Z(
        n1681) );
  HS65_LL_OAI21X3 U14810 ( .A(n3054), .B(n3225), .C(n4080), .Z(n4106) );
  HS65_LL_NAND4ABX3 U14811 ( .A(n6845), .B(n6846), .C(n6847), .D(n6848), .Z(
        n6320) );
  HS65_LL_NOR3AX2 U14812 ( .A(n6853), .B(n6854), .C(n6855), .Z(n6847) );
  HS65_LL_OAI212X5 U14813 ( .A(n6856), .B(n6857), .C(n6476), .D(n6047), .E(
        n6858), .Z(n6846) );
  HS65_LL_NOR4ABX2 U14814 ( .A(n6849), .B(n6850), .C(n6851), .D(n6852), .Z(
        n6848) );
  HS65_LL_NAND4ABX3 U14815 ( .A(n5253), .B(n5254), .C(n5255), .D(n5256), .Z(
        n4740) );
  HS65_LL_NOR3AX2 U14816 ( .A(n5261), .B(n5262), .C(n5263), .Z(n5255) );
  HS65_LL_OAI212X5 U14817 ( .A(n5264), .B(n5265), .C(n4883), .D(n4454), .E(
        n5266), .Z(n5254) );
  HS65_LL_NOR4ABX2 U14818 ( .A(n5257), .B(n5258), .C(n5259), .D(n5260), .Z(
        n5256) );
  HS65_LL_IVX9 U14819 ( .A(n7847), .Z(n378) );
  HS65_LL_IVX9 U14820 ( .A(n2333), .Z(n902) );
  HS65_LL_IVX9 U14821 ( .A(n1581), .Z(n820) );
  HS65_LL_IVX9 U14822 ( .A(n1205), .Z(n861) );
  HS65_LL_IVX9 U14823 ( .A(n1957), .Z(n779) );
  HS65_LL_IVX9 U14824 ( .A(n7947), .Z(n317) );
  HS65_LL_IVX9 U14825 ( .A(n2361), .Z(n911) );
  HS65_LL_IVX9 U14826 ( .A(n1609), .Z(n829) );
  HS65_LL_IVX9 U14827 ( .A(n1233), .Z(n870) );
  HS65_LL_IVX9 U14828 ( .A(n1985), .Z(n788) );
  HS65_LL_IVX9 U14829 ( .A(n2888), .Z(n638) );
  HS65_LL_IVX9 U14830 ( .A(n3380), .Z(n412) );
  HS65_LL_NOR2X6 U14831 ( .A(n3158), .B(n2972), .Z(n3710) );
  HS65_LL_NOR2X6 U14832 ( .A(n3185), .B(n2997), .Z(n3825) );
  HS65_LL_NOR2X6 U14833 ( .A(n2958), .B(n2859), .Z(n3469) );
  HS65_LL_NAND2X7 U14834 ( .A(n1895), .B(n1862), .Z(n2038) );
  HS65_LL_NAND2X7 U14835 ( .A(n1143), .B(n1110), .Z(n1286) );
  HS65_LL_NOR2X6 U14836 ( .A(n7750), .B(n7980), .Z(n8113) );
  HS65_LL_NOR2X6 U14837 ( .A(n7768), .B(n8048), .Z(n8346) );
  HS65_LL_NOR2X6 U14838 ( .A(n5267), .B(n4748), .Z(n4759) );
  HS65_LL_NOR2X6 U14839 ( .A(n5382), .B(n4774), .Z(n4786) );
  HS65_LL_NOR2X6 U14840 ( .A(n6974), .B(n6367), .Z(n6379) );
  HS65_LL_NOR2X6 U14841 ( .A(n6859), .B(n6328), .Z(n6340) );
  HS65_LL_IVX9 U14842 ( .A(n3067), .Z(n196) );
  HS65_LL_NAND2X7 U14843 ( .A(n1143), .B(n1233), .Z(n1301) );
  HS65_LL_NAND2X7 U14844 ( .A(n1895), .B(n1985), .Z(n2053) );
  HS65_LL_NAND2X7 U14845 ( .A(n4589), .B(n250), .Z(n4753) );
  HS65_LL_NAND2X7 U14846 ( .A(n6182), .B(n91), .Z(n6334) );
  HS65_LL_IVX9 U14847 ( .A(n2931), .Z(n195) );
  HS65_LL_NOR2X6 U14848 ( .A(n3807), .B(n3846), .Z(n3815) );
  HS65_LL_IVX9 U14849 ( .A(n8155), .Z(n587) );
  HS65_LL_IVX9 U14850 ( .A(n8178), .Z(n107) );
  HS65_LL_IVX9 U14851 ( .A(n3096), .Z(n199) );
  HS65_LL_NOR2X6 U14852 ( .A(n4477), .B(n5507), .Z(n4573) );
  HS65_LL_NOR2X6 U14853 ( .A(n6070), .B(n7099), .Z(n6166) );
  HS65_LL_IVX9 U14854 ( .A(n1537), .Z(n828) );
  HS65_LL_NOR2X6 U14855 ( .A(n7686), .B(n7623), .Z(n8418) );
  HS65_LL_NOR2X6 U14856 ( .A(n7724), .B(n7663), .Z(n8470) );
  HS65_LL_NAND2X7 U14857 ( .A(n264), .B(n4589), .Z(n5321) );
  HS65_LL_NAND2X7 U14858 ( .A(n481), .B(n4606), .Z(n5436) );
  HS65_LL_NAND2X7 U14859 ( .A(n78), .B(n6182), .Z(n6913) );
  HS65_LL_NAND2X7 U14860 ( .A(n306), .B(n6199), .Z(n7028) );
  HS65_LL_NOR2X6 U14861 ( .A(n1743), .B(n1695), .Z(n1665) );
  HS65_LL_NOR2X6 U14862 ( .A(n2495), .B(n2447), .Z(n2417) );
  HS65_LL_IVX9 U14863 ( .A(n2289), .Z(n910) );
  HS65_LL_NOR2X6 U14864 ( .A(n2119), .B(n2071), .Z(n2041) );
  HS65_LL_NOR2X6 U14865 ( .A(n1367), .B(n1319), .Z(n1289) );
  HS65_LL_IVX9 U14866 ( .A(n1913), .Z(n787) );
  HS65_LL_IVX9 U14867 ( .A(n1161), .Z(n869) );
  HS65_LL_NOR2X6 U14868 ( .A(n2308), .B(n2257), .Z(n2367) );
  HS65_LL_NOR2X6 U14869 ( .A(n1556), .B(n1505), .Z(n1615) );
  HS65_LL_NOR2X6 U14870 ( .A(n1932), .B(n1881), .Z(n1991) );
  HS65_LL_NOR2X6 U14871 ( .A(n1180), .B(n1129), .Z(n1239) );
  HS65_LL_OAI21X3 U14872 ( .A(n7882), .B(n7713), .C(n7733), .Z(n7881) );
  HS65_LL_OAI21X3 U14873 ( .A(n7783), .B(n7675), .C(n7695), .Z(n7782) );
  HS65_LL_IVX9 U14874 ( .A(n4923), .Z(n235) );
  HS65_LL_IVX9 U14875 ( .A(n6569), .Z(n277) );
  HS65_LL_IVX9 U14876 ( .A(n6516), .Z(n66) );
  HS65_LL_IVX9 U14877 ( .A(n4976), .Z(n452) );
  HS65_LL_NOR2X6 U14878 ( .A(n8058), .B(n8540), .Z(n8511) );
  HS65_LL_NOR2X6 U14879 ( .A(n3185), .B(n2845), .Z(n3386) );
  HS65_LL_NOR2X6 U14880 ( .A(n3158), .B(n2875), .Z(n3332) );
  HS65_LL_NOR2X6 U14881 ( .A(n8028), .B(n7942), .Z(n8500) );
  HS65_LL_NAND3X5 U14882 ( .A(n1168), .B(n1199), .C(n1155), .Z(n1419) );
  HS65_LL_IVX9 U14883 ( .A(n3197), .Z(n416) );
  HS65_LL_IVX9 U14884 ( .A(n4670), .Z(n11) );
  HS65_LL_IVX9 U14885 ( .A(n6263), .Z(n533) );
  HS65_LL_NAND2X7 U14886 ( .A(n4589), .B(n265), .Z(n4925) );
  HS65_LL_NAND2X7 U14887 ( .A(n6182), .B(n79), .Z(n6518) );
  HS65_LL_NOR2X6 U14888 ( .A(n6515), .B(n6327), .Z(n6922) );
  HS65_LL_NOR2X6 U14889 ( .A(n4922), .B(n4747), .Z(n5330) );
  HS65_LL_NOR2X6 U14890 ( .A(n4975), .B(n4773), .Z(n5445) );
  HS65_LL_NOR2X6 U14891 ( .A(n6568), .B(n6366), .Z(n7037) );
  HS65_LL_NOR2X6 U14892 ( .A(n1985), .B(n1863), .Z(n2002) );
  HS65_LL_NAND2X7 U14893 ( .A(n473), .B(n4606), .Z(n5373) );
  HS65_LL_NAND2X7 U14894 ( .A(n256), .B(n4589), .Z(n5258) );
  HS65_LL_NAND2X7 U14895 ( .A(n74), .B(n6182), .Z(n6850) );
  HS65_LL_NAND2X7 U14896 ( .A(n298), .B(n6199), .Z(n6965) );
  HS65_LL_NOR2X6 U14897 ( .A(n2958), .B(n2940), .Z(n3103) );
  HS65_LL_NOR4ABX2 U14898 ( .A(n5521), .B(n5529), .C(n4452), .D(n5590), .Z(
        n5585) );
  HS65_LL_OAI212X5 U14899 ( .A(n5533), .B(n4455), .C(n5591), .D(n4460), .E(
        n5592), .Z(n5590) );
  HS65_LL_NOR4ABX2 U14900 ( .A(n7113), .B(n7121), .C(n6045), .D(n7182), .Z(
        n7177) );
  HS65_LL_OAI212X5 U14901 ( .A(n7125), .B(n6048), .C(n7183), .D(n6053), .E(
        n7184), .Z(n7182) );
  HS65_LL_IVX9 U14902 ( .A(n6328), .Z(n91) );
  HS65_LL_NOR2X6 U14903 ( .A(n2361), .B(n2239), .Z(n2378) );
  HS65_LL_NOR2X6 U14904 ( .A(n1233), .B(n1111), .Z(n1250) );
  HS65_LL_NOR2X6 U14905 ( .A(n1609), .B(n1487), .Z(n1626) );
  HS65_LL_NAND2X7 U14906 ( .A(n252), .B(n4589), .Z(n5276) );
  HS65_LL_NAND2X7 U14907 ( .A(n89), .B(n6182), .Z(n6868) );
  HS65_LL_NOR4ABX2 U14908 ( .A(n3937), .B(n3938), .C(n3939), .D(n3940), .Z(
        n3932) );
  HS65_LL_OAI212X5 U14909 ( .A(n3293), .B(n3342), .C(n3158), .D(n2884), .E(
        n2878), .Z(n3939) );
  HS65_LL_NOR2X6 U14910 ( .A(n3157), .B(n2888), .Z(n3699) );
  HS65_LL_NOR4ABX2 U14911 ( .A(n3892), .B(n3893), .C(n3894), .D(n3895), .Z(
        n3887) );
  HS65_LL_OAI212X5 U14912 ( .A(n3061), .B(n3114), .C(n2958), .D(n2956), .E(
        n3896), .Z(n3895) );
  HS65_LL_NOR2X6 U14913 ( .A(n3183), .B(n2836), .Z(n3814) );
  HS65_LL_NAND2X7 U14914 ( .A(n609), .B(n7699), .Z(n8696) );
  HS65_LL_NAND2X7 U14915 ( .A(n129), .B(n7737), .Z(n8786) );
  HS65_LL_NOR2X6 U14916 ( .A(n8510), .B(n8039), .Z(n8353) );
  HS65_LL_NOR2X6 U14917 ( .A(n8207), .B(n7971), .Z(n8077) );
  HS65_LL_NOR4ABX2 U14918 ( .A(n3937), .B(n4001), .C(n2880), .D(n4002), .Z(
        n3997) );
  HS65_LL_OA212X4 U14919 ( .A(n2884), .B(n3141), .C(n3692), .D(n2888), .E(
        n3947), .Z(n4001) );
  HS65_LL_NOR4ABX2 U14920 ( .A(n7854), .B(n7855), .C(n7856), .D(n7857), .Z(
        n7843) );
  HS65_LL_OA212X4 U14921 ( .A(n7858), .B(n7859), .C(n7860), .D(n7861), .E(
        n7862), .Z(n7854) );
  HS65_LL_NAND4ABX3 U14922 ( .A(n1973), .B(n1974), .C(n1975), .D(n1976), .Z(
        n1893) );
  HS65_LL_OAI222X2 U14923 ( .A(n1863), .B(n1897), .C(n1932), .D(n1985), .E(
        n1881), .F(n1861), .Z(n1974) );
  HS65_LL_NOR4ABX2 U14924 ( .A(n1981), .B(n1982), .C(n1983), .D(n1984), .Z(
        n1975) );
  HS65_LL_NOR4ABX2 U14925 ( .A(n1977), .B(n1978), .C(n1979), .D(n1980), .Z(
        n1976) );
  HS65_LL_NAND4ABX3 U14926 ( .A(n2349), .B(n2350), .C(n2351), .D(n2352), .Z(
        n2269) );
  HS65_LL_OAI222X2 U14927 ( .A(n2239), .B(n2273), .C(n2308), .D(n2361), .E(
        n2257), .F(n2237), .Z(n2350) );
  HS65_LL_NOR4ABX2 U14928 ( .A(n2357), .B(n2358), .C(n2359), .D(n2360), .Z(
        n2351) );
  HS65_LL_NOR4ABX2 U14929 ( .A(n2353), .B(n2354), .C(n2355), .D(n2356), .Z(
        n2352) );
  HS65_LL_NAND4ABX3 U14930 ( .A(n1221), .B(n1222), .C(n1223), .D(n1224), .Z(
        n1141) );
  HS65_LL_OAI222X2 U14931 ( .A(n1111), .B(n1145), .C(n1180), .D(n1233), .E(
        n1129), .F(n1109), .Z(n1222) );
  HS65_LL_NOR4ABX2 U14932 ( .A(n1229), .B(n1230), .C(n1231), .D(n1232), .Z(
        n1223) );
  HS65_LL_NOR4ABX2 U14933 ( .A(n1225), .B(n1226), .C(n1227), .D(n1228), .Z(
        n1224) );
  HS65_LL_NAND4ABX3 U14934 ( .A(n1597), .B(n1598), .C(n1599), .D(n1600), .Z(
        n1517) );
  HS65_LL_OAI222X2 U14935 ( .A(n1487), .B(n1521), .C(n1556), .D(n1609), .E(
        n1505), .F(n1485), .Z(n1598) );
  HS65_LL_NOR4ABX2 U14936 ( .A(n1605), .B(n1606), .C(n1607), .D(n1608), .Z(
        n1599) );
  HS65_LL_NOR4ABX2 U14937 ( .A(n1601), .B(n1602), .C(n1603), .D(n1604), .Z(
        n1600) );
  HS65_LL_NAND4ABX3 U14938 ( .A(n3314), .B(n3315), .C(n3316), .D(n3317), .Z(
        n2979) );
  HS65_LL_OAI222X2 U14939 ( .A(n2883), .B(n2969), .C(n3158), .D(n3326), .E(
        n2875), .F(n2881), .Z(n3315) );
  HS65_LL_NOR4ABX2 U14940 ( .A(n3318), .B(n3319), .C(n3320), .D(n3321), .Z(
        n3317) );
  HS65_LL_NAND3AX6 U14941 ( .A(n3327), .B(n3328), .C(n3329), .Z(n3314) );
  HS65_LL_NOR2X6 U14942 ( .A(n6159), .B(n7093), .Z(n6595) );
  HS65_LL_NOR2X6 U14943 ( .A(n4566), .B(n5501), .Z(n5002) );
  HS65_LL_NOR4ABX2 U14944 ( .A(n7626), .B(n7627), .C(n7628), .D(n7629), .Z(
        n7615) );
  HS65_LL_OA212X4 U14945 ( .A(n7630), .B(n7631), .C(n7632), .D(n7633), .E(
        n7634), .Z(n7627) );
  HS65_LL_IVX9 U14946 ( .A(n4478), .Z(n23) );
  HS65_LL_IVX9 U14947 ( .A(n6071), .Z(n545) );
  HS65_LL_IVX9 U14948 ( .A(n4454), .Z(n233) );
  HS65_LL_IVX9 U14949 ( .A(n4493), .Z(n450) );
  HS65_LL_IVX9 U14950 ( .A(n6047), .Z(n64) );
  HS65_LL_IVX9 U14951 ( .A(n6086), .Z(n275) );
  HS65_LL_IVX9 U14952 ( .A(n6127), .Z(n502) );
  HS65_LL_NAND2X7 U14953 ( .A(n4589), .B(n257), .Z(n4918) );
  HS65_LL_NAND2X7 U14954 ( .A(n6182), .B(n76), .Z(n6511) );
  HS65_LL_NOR3AX2 U14955 ( .A(n8621), .B(n8885), .C(n8857), .Z(n8879) );
  HS65_LL_OAI21X3 U14956 ( .A(n8033), .B(n8049), .C(n8869), .Z(n8885) );
  HS65_LL_NOR3AX2 U14957 ( .A(n8636), .B(n8945), .C(n8644), .Z(n8939) );
  HS65_LL_OAI21X3 U14958 ( .A(n7965), .B(n7981), .C(n8491), .Z(n8945) );
  HS65_LL_NAND4ABX3 U14959 ( .A(n2131), .B(n2132), .C(n2133), .D(n2134), .Z(
        n2129) );
  HS65_LL_OA212X4 U14960 ( .A(n2121), .B(n1951), .C(n1864), .D(n1932), .E(
        n1878), .Z(n2134) );
  HS65_LL_NAND4ABX3 U14961 ( .A(n1379), .B(n1380), .C(n1381), .D(n1382), .Z(
        n1377) );
  HS65_LL_OA212X4 U14962 ( .A(n1369), .B(n1199), .C(n1112), .D(n1180), .E(
        n1126), .Z(n1382) );
  HS65_LL_NAND4ABX3 U14963 ( .A(n2507), .B(n2508), .C(n2509), .D(n2510), .Z(
        n2505) );
  HS65_LL_OA212X4 U14964 ( .A(n2497), .B(n2327), .C(n2240), .D(n2308), .E(
        n2254), .Z(n2510) );
  HS65_LL_NAND4ABX3 U14965 ( .A(n1755), .B(n1756), .C(n1757), .D(n1758), .Z(
        n1753) );
  HS65_LL_OA212X4 U14966 ( .A(n1745), .B(n1575), .C(n1488), .D(n1556), .E(
        n1502), .Z(n1758) );
  HS65_LL_NOR4ABX2 U14967 ( .A(n9072), .B(n8798), .C(n8436), .D(n8815), .Z(
        n9069) );
  HS65_LL_OAI21X3 U14968 ( .A(n98), .B(n7737), .C(n136), .Z(n9072) );
  HS65_LL_NOR4ABX2 U14969 ( .A(n9014), .B(n8708), .C(n8384), .D(n8725), .Z(
        n9011) );
  HS65_LL_OAI21X3 U14970 ( .A(n578), .B(n7699), .C(n616), .Z(n9014) );
  HS65_LL_NOR4ABX2 U14971 ( .A(n5898), .B(n5463), .C(n5420), .D(n4959), .Z(
        n5895) );
  HS65_LL_OAI21X3 U14972 ( .A(n461), .B(n4606), .C(n476), .Z(n5898) );
  HS65_LL_NOR4ABX2 U14973 ( .A(n5839), .B(n5348), .C(n5305), .D(n4906), .Z(
        n5836) );
  HS65_LL_OAI21X3 U14974 ( .A(n244), .B(n4589), .C(n259), .Z(n5839) );
  HS65_LL_NOR4ABX2 U14975 ( .A(n7490), .B(n7055), .C(n7012), .D(n6552), .Z(
        n7487) );
  HS65_LL_OAI21X3 U14976 ( .A(n286), .B(n6199), .C(n301), .Z(n7490) );
  HS65_LL_NOR4ABX2 U14977 ( .A(n5799), .B(n5233), .C(n5189), .D(n4831), .Z(
        n5796) );
  HS65_LL_OAI21X3 U14978 ( .A(n670), .B(n4521), .C(n685), .Z(n5799) );
  HS65_LL_NOR4ABX2 U14979 ( .A(n7391), .B(n6825), .C(n6781), .D(n6424), .Z(
        n7388) );
  HS65_LL_OAI21X3 U14980 ( .A(n494), .B(n6114), .C(n509), .Z(n7391) );
  HS65_LL_NOR4ABX2 U14981 ( .A(n7431), .B(n6940), .C(n6897), .D(n6499), .Z(
        n7428) );
  HS65_LL_OAI21X3 U14982 ( .A(n55), .B(n6182), .C(n77), .Z(n7431) );
  HS65_LL_NAND2X7 U14983 ( .A(n563), .B(n6074), .Z(n6270) );
  HS65_LL_NAND2X7 U14984 ( .A(n41), .B(n4481), .Z(n4677) );
  HS65_LL_IVX9 U14985 ( .A(n5267), .Z(n238) );
  HS65_LL_IVX9 U14986 ( .A(n6974), .Z(n280) );
  HS65_LL_IVX9 U14987 ( .A(n6859), .Z(n60) );
  HS65_LL_NAND4ABX3 U14988 ( .A(n1124), .B(n1125), .C(n1126), .D(n1127), .Z(
        n1106) );
  HS65_LL_AOI212X4 U14989 ( .A(n866), .B(n845), .C(n874), .D(n850), .E(n1128), 
        .Z(n1127) );
  HS65_LL_OAI21X3 U14990 ( .A(n1129), .B(n1130), .C(n1131), .Z(n1128) );
  HS65_LL_NAND4ABX3 U14991 ( .A(n1876), .B(n1877), .C(n1878), .D(n1879), .Z(
        n1858) );
  HS65_LL_AOI212X4 U14992 ( .A(n784), .B(n763), .C(n792), .D(n768), .E(n1880), 
        .Z(n1879) );
  HS65_LL_OAI21X3 U14993 ( .A(n1881), .B(n1882), .C(n1883), .Z(n1880) );
  HS65_LL_NAND4ABX3 U14994 ( .A(n2268), .B(n2299), .C(n2334), .D(n2335), .Z(
        n2322) );
  HS65_LL_AOI212X4 U14995 ( .A(n901), .B(n887), .C(n894), .D(n902), .E(n2336), 
        .Z(n2335) );
  HS65_LL_OAI21X3 U14996 ( .A(n2257), .B(n2246), .C(n2337), .Z(n2336) );
  HS65_LL_NAND4ABX3 U14997 ( .A(n1892), .B(n1923), .C(n1958), .D(n1959), .Z(
        n1946) );
  HS65_LL_AOI212X4 U14998 ( .A(n778), .B(n764), .C(n771), .D(n779), .E(n1960), 
        .Z(n1959) );
  HS65_LL_OAI21X3 U14999 ( .A(n1881), .B(n1870), .C(n1961), .Z(n1960) );
  HS65_LL_NAND4ABX3 U15000 ( .A(n1140), .B(n1171), .C(n1206), .D(n1207), .Z(
        n1194) );
  HS65_LL_AOI212X4 U15001 ( .A(n860), .B(n846), .C(n853), .D(n861), .E(n1208), 
        .Z(n1207) );
  HS65_LL_OAI21X3 U15002 ( .A(n1129), .B(n1118), .C(n1209), .Z(n1208) );
  HS65_LL_NAND4ABX3 U15003 ( .A(n1516), .B(n1547), .C(n1582), .D(n1583), .Z(
        n1570) );
  HS65_LL_AOI212X4 U15004 ( .A(n819), .B(n805), .C(n812), .D(n820), .E(n1584), 
        .Z(n1583) );
  HS65_LL_OAI21X3 U15005 ( .A(n1505), .B(n1494), .C(n1585), .Z(n1584) );
  HS65_LL_NAND4ABX3 U15006 ( .A(n1500), .B(n1501), .C(n1502), .D(n1503), .Z(
        n1482) );
  HS65_LL_AOI212X4 U15007 ( .A(n825), .B(n804), .C(n833), .D(n809), .E(n1504), 
        .Z(n1503) );
  HS65_LL_OAI21X3 U15008 ( .A(n1505), .B(n1506), .C(n1507), .Z(n1504) );
  HS65_LL_NAND4ABX3 U15009 ( .A(n2252), .B(n2253), .C(n2254), .D(n2255), .Z(
        n2234) );
  HS65_LL_AOI212X4 U15010 ( .A(n907), .B(n886), .C(n915), .D(n891), .E(n2256), 
        .Z(n2255) );
  HS65_LL_OAI21X3 U15011 ( .A(n2257), .B(n2258), .C(n2259), .Z(n2256) );
  HS65_LL_NAND2X7 U15012 ( .A(n309), .B(n6199), .Z(n6537) );
  HS65_LL_NAND2X7 U15013 ( .A(n81), .B(n6182), .Z(n6484) );
  HS65_LL_NAND2X7 U15014 ( .A(n267), .B(n4589), .Z(n4891) );
  HS65_LL_NAND2X7 U15015 ( .A(n484), .B(n4606), .Z(n4944) );
  HS65_LL_NAND2X7 U15016 ( .A(n520), .B(n6114), .Z(n6409) );
  HS65_LL_NAND2X7 U15017 ( .A(n696), .B(n4521), .Z(n4816) );
  HS65_LL_OAI212X5 U15018 ( .A(n1629), .B(n1506), .C(n1532), .D(n1494), .E(
        n1630), .Z(n1619) );
  HS65_LL_NOR2X6 U15019 ( .A(n831), .B(n820), .Z(n1629) );
  HS65_LL_OAI21X3 U15020 ( .A(n833), .B(n827), .C(n807), .Z(n1630) );
  HS65_LL_OAI212X5 U15021 ( .A(n2381), .B(n2258), .C(n2284), .D(n2246), .E(
        n2382), .Z(n2371) );
  HS65_LL_NOR2X6 U15022 ( .A(n913), .B(n902), .Z(n2381) );
  HS65_LL_OAI21X3 U15023 ( .A(n915), .B(n909), .C(n889), .Z(n2382) );
  HS65_LL_NOR4ABX2 U15024 ( .A(n5737), .B(n5097), .C(n5067), .D(n4693), .Z(
        n5734) );
  HS65_LL_OAI21X3 U15025 ( .A(n15), .B(n4481), .C(n30), .Z(n5737) );
  HS65_LL_NOR4ABX2 U15026 ( .A(n7329), .B(n6690), .C(n6660), .D(n6286), .Z(
        n7326) );
  HS65_LL_OAI21X3 U15027 ( .A(n537), .B(n6074), .C(n552), .Z(n7329) );
  HS65_LL_IVX9 U15028 ( .A(n4882), .Z(n232) );
  HS65_LL_IVX9 U15029 ( .A(n4994), .Z(n449) );
  HS65_LL_IVX9 U15030 ( .A(n6475), .Z(n65) );
  HS65_LL_IVX9 U15031 ( .A(n6587), .Z(n274) );
  HS65_LL_OAI212X5 U15032 ( .A(n2535), .B(n2244), .C(n2445), .D(n2271), .E(
        n2536), .Z(n2534) );
  HS65_LL_NOR3X4 U15033 ( .A(n882), .B(n891), .C(n884), .Z(n2535) );
  HS65_LL_OAI21X3 U15034 ( .A(n907), .B(n914), .C(n896), .Z(n2536) );
  HS65_LL_OAI212X5 U15035 ( .A(n7189), .B(n6053), .C(n6186), .D(n6857), .E(
        n7190), .Z(n7188) );
  HS65_LL_NOR3X4 U15036 ( .A(n86), .B(n91), .C(n90), .Z(n7189) );
  HS65_LL_OAI21X3 U15037 ( .A(n63), .B(n56), .C(n79), .Z(n7190) );
  HS65_LL_OAI212X5 U15038 ( .A(n4007), .B(n2888), .C(n3343), .D(n2981), .E(
        n4008), .Z(n4006) );
  HS65_LL_NOR3X4 U15039 ( .A(n656), .B(n648), .C(n644), .Z(n4007) );
  HS65_LL_OAI21X3 U15040 ( .A(n631), .B(n635), .C(n660), .Z(n4008) );
  HS65_LL_AOI12X2 U15041 ( .A(n839), .B(n1159), .C(n1160), .Z(n1158) );
  HS65_LL_AOI12X2 U15042 ( .A(n1161), .B(n1162), .C(n1163), .Z(n1160) );
  HS65_LL_OAI21X3 U15043 ( .A(n8150), .B(n7831), .C(n8727), .Z(n9009) );
  HS65_LL_OAI21X3 U15044 ( .A(n8173), .B(n7870), .C(n8817), .Z(n9067) );
  HS65_LL_OAI21X3 U15045 ( .A(n4994), .B(n4495), .C(n5458), .Z(n5919) );
  HS65_LL_OAI21X3 U15046 ( .A(n6587), .B(n6088), .C(n7050), .Z(n7511) );
  HS65_LL_OAI21X3 U15047 ( .A(n4882), .B(n4456), .C(n5343), .Z(n5860) );
  HS65_LL_OAI21X3 U15048 ( .A(n6475), .B(n6049), .C(n6935), .Z(n7452) );
  HS65_LL_OAI21X3 U15049 ( .A(n4868), .B(n4848), .C(n5228), .Z(n5788) );
  HS65_LL_OAI21X3 U15050 ( .A(n6461), .B(n6441), .C(n6820), .Z(n7380) );
  HS65_LL_NAND2X7 U15051 ( .A(n7699), .B(n610), .Z(n8408) );
  HS65_LL_NAND2X7 U15052 ( .A(n7737), .B(n130), .Z(n8460) );
  HS65_LL_OAI21X3 U15053 ( .A(n6260), .B(n6302), .C(n6685), .Z(n7318) );
  HS65_LL_OAI21X3 U15054 ( .A(n4667), .B(n4709), .C(n5092), .Z(n5726) );
  HS65_LL_OAI212X5 U15055 ( .A(n8687), .B(n7822), .C(n8421), .D(n7806), .E(
        n8688), .Z(n8679) );
  HS65_LL_NOR2X6 U15056 ( .A(n576), .B(n8666), .Z(n8687) );
  HS65_LL_OAI212X5 U15057 ( .A(n8777), .B(n7920), .C(n8473), .D(n7869), .E(
        n8778), .Z(n8769) );
  HS65_LL_NOR2X6 U15058 ( .A(n96), .B(n8756), .Z(n8777) );
  HS65_LL_OAI212X5 U15059 ( .A(n3729), .B(n3343), .C(n2970), .D(n2882), .E(
        n3730), .Z(n3719) );
  HS65_LL_NOR2X6 U15060 ( .A(n634), .B(n3660), .Z(n3729) );
  HS65_LL_OAI212X5 U15061 ( .A(n8252), .B(n7993), .C(n7848), .D(n7851), .E(
        n8253), .Z(n8242) );
  HS65_LL_NOR2X6 U15062 ( .A(n368), .B(n8195), .Z(n8252) );
  HS65_LL_MX41X7 U15063 ( .D0(n585), .S0(n602), .D1(n616), .S1(n593), .D2(n605), .S2(n7699), .D3(n588), .S3(n612), .Z(n8743) );
  HS65_LL_CB4I1X9 U15064 ( .A(n2146), .B(n1921), .C(n2071), .D(n2122), .Z(
        n2170) );
  HS65_LL_OAI212X5 U15065 ( .A(n1368), .B(n1129), .C(n1146), .D(n1233), .E(
        n1418), .Z(n1416) );
  HS65_LL_CB4I1X9 U15066 ( .A(n1394), .B(n1169), .C(n1319), .D(n1370), .Z(
        n1418) );
  HS65_LL_CB4I1X9 U15067 ( .A(n2522), .B(n2297), .C(n2447), .D(n2498), .Z(
        n2546) );
  HS65_LL_CB4I1X9 U15068 ( .A(n1770), .B(n1545), .C(n1695), .D(n1746), .Z(
        n1794) );
  HS65_LL_AND2X4 U15069 ( .A(n7699), .B(n604), .Z(n8151) );
  HS65_LL_OA12X9 U15070 ( .A(n8510), .B(n7949), .C(n8586), .Z(n8585) );
  HS65_LL_AND2X4 U15071 ( .A(n4589), .B(n263), .Z(n4751) );
  HS65_LL_AND2X4 U15072 ( .A(n4606), .B(n480), .Z(n4778) );
  HS65_LL_AND2X4 U15073 ( .A(n6199), .B(n305), .Z(n6371) );
  HS65_LL_AND2X4 U15074 ( .A(n6182), .B(n86), .Z(n6332) );
  HS65_LL_NOR4ABX2 U15075 ( .A(n8023), .B(n8024), .C(n8025), .D(n8026), .Z(
        n3003) );
  HS65_LL_NAND4ABX3 U15076 ( .A(n8035), .B(n8036), .C(n8037), .D(n8038), .Z(
        n8025) );
  HS65_LL_OAI212X5 U15077 ( .A(n8027), .B(n8028), .C(n8029), .D(n7952), .E(
        n8030), .Z(n8026) );
  HS65_LL_AOI212X4 U15078 ( .A(n349), .B(n322), .C(n333), .D(n356), .E(n8040), 
        .Z(n8024) );
  HS65_LL_NOR4ABX2 U15079 ( .A(n8477), .B(n8478), .C(n8479), .D(n8480), .Z(
        n2752) );
  HS65_LL_CB4I6X9 U15080 ( .A(n393), .B(n398), .C(n378), .D(n8273), .Z(n8479)
         );
  HS65_LL_CBI4I1X5 U15081 ( .A(n8481), .B(n7751), .C(n7850), .D(n8482), .Z(
        n8480) );
  HS65_LL_AOI212X4 U15082 ( .A(n371), .B(n399), .C(n373), .D(n8492), .E(n8493), 
        .Z(n8477) );
  HS65_LL_NOR4ABX2 U15083 ( .A(n5466), .B(n5467), .C(n5468), .D(n5469), .Z(
        n2768) );
  HS65_LL_CBI4I1X5 U15084 ( .A(n4572), .B(n4709), .C(n4710), .D(n5046), .Z(
        n5468) );
  HS65_LL_CBI4I1X5 U15085 ( .A(n5470), .B(n4712), .C(n4477), .D(n5471), .Z(
        n5469) );
  HS65_LL_AOI212X4 U15086 ( .A(n18), .B(n37), .C(n19), .D(n5478), .E(n5479), 
        .Z(n5466) );
  HS65_LL_NOR4ABX2 U15087 ( .A(n7058), .B(n7059), .C(n7060), .D(n7061), .Z(
        n2760) );
  HS65_LL_CBI4I1X5 U15088 ( .A(n6165), .B(n6302), .C(n6303), .D(n6639), .Z(
        n7060) );
  HS65_LL_CBI4I1X5 U15089 ( .A(n7062), .B(n6305), .C(n6070), .D(n7063), .Z(
        n7061) );
  HS65_LL_AOI212X4 U15090 ( .A(n540), .B(n559), .C(n541), .D(n7070), .E(n7071), 
        .Z(n7058) );
  HS65_LL_IVX9 U15091 ( .A(n3047), .Z(n150) );
  HS65_LL_NOR4ABX2 U15092 ( .A(n2921), .B(n2922), .C(n2923), .D(n2924), .Z(
        n2644) );
  HS65_LL_NAND4ABX3 U15093 ( .A(n2934), .B(n2935), .C(n2936), .D(n2937), .Z(
        n2923) );
  HS65_LL_OAI212X5 U15094 ( .A(n2925), .B(n2926), .C(n2927), .D(n2860), .E(
        n2928), .Z(n2924) );
  HS65_LL_AOI212X4 U15095 ( .A(n188), .B(n213), .C(n192), .D(n219), .E(n2941), 
        .Z(n2922) );
  HS65_LL_NOR4ABX2 U15096 ( .A(n3123), .B(n3124), .C(n3125), .D(n3126), .Z(
        n2634) );
  HS65_LL_NAND4ABX3 U15097 ( .A(n3136), .B(n3137), .C(n3138), .D(n3139), .Z(
        n3125) );
  HS65_LL_OAI212X5 U15098 ( .A(n3127), .B(n3128), .C(n3129), .D(n2882), .E(
        n3130), .Z(n3126) );
  HS65_LL_AOI212X4 U15099 ( .A(n638), .B(n656), .C(n633), .D(n651), .E(n3142), 
        .Z(n3124) );
  HS65_LL_NAND4ABX3 U15100 ( .A(n8062), .B(n8063), .C(n8064), .D(n8065), .Z(
        n2754) );
  HS65_LL_NAND4ABX3 U15101 ( .A(n8119), .B(n8120), .C(n8121), .D(n8122), .Z(
        n8062) );
  HS65_LL_OAI212X5 U15102 ( .A(n8116), .B(n7861), .C(n7752), .D(n8117), .E(
        n8118), .Z(n8063) );
  HS65_LL_AOI212X4 U15103 ( .A(n373), .B(n388), .C(n377), .D(n383), .E(n8066), 
        .Z(n8065) );
  HS65_LL_NAND4ABX3 U15104 ( .A(n8422), .B(n8423), .C(n8424), .D(n8425), .Z(
        n2802) );
  HS65_LL_NAND4ABX3 U15105 ( .A(n8469), .B(n8470), .C(n8471), .D(n8472), .Z(
        n8422) );
  HS65_LL_OAI212X5 U15106 ( .A(n8467), .B(n7650), .C(n7715), .D(n7657), .E(
        n8468), .Z(n8423) );
  HS65_LL_AOI212X4 U15107 ( .A(n112), .B(n128), .C(n108), .D(n122), .E(n8426), 
        .Z(n8425) );
  HS65_LL_NAND4ABX3 U15108 ( .A(n6207), .B(n6208), .C(n6209), .D(n6210), .Z(
        n3206) );
  HS65_LL_NAND4ABX3 U15109 ( .A(n6243), .B(n6244), .C(n6245), .D(n6246), .Z(
        n6207) );
  HS65_LL_OAI212X5 U15110 ( .A(n6235), .B(n6236), .C(n6127), .D(n6237), .E(
        n6238), .Z(n6208) );
  HS65_LL_AOI212X4 U15111 ( .A(n489), .B(n513), .C(n509), .D(n493), .E(n6211), 
        .Z(n6210) );
  HS65_LL_NAND4ABX3 U15112 ( .A(n4614), .B(n4615), .C(n4616), .D(n4617), .Z(
        n3214) );
  HS65_LL_NAND4ABX3 U15113 ( .A(n4650), .B(n4651), .C(n4652), .D(n4653), .Z(
        n4614) );
  HS65_LL_OAI212X5 U15114 ( .A(n4642), .B(n4643), .C(n4534), .D(n4644), .E(
        n4645), .Z(n4615) );
  HS65_LL_AOI212X4 U15115 ( .A(n665), .B(n689), .C(n685), .D(n669), .E(n4618), 
        .Z(n4617) );
  HS65_LL_NAND4ABX3 U15116 ( .A(n6315), .B(n6316), .C(n6317), .D(n6318), .Z(
        n2787) );
  HS65_LL_NAND4ABX3 U15117 ( .A(n6350), .B(n6351), .C(n6352), .D(n6353), .Z(
        n6315) );
  HS65_LL_OAI212X5 U15118 ( .A(n6342), .B(n6343), .C(n6047), .D(n6344), .E(
        n6345), .Z(n6316) );
  HS65_LL_AOI212X4 U15119 ( .A(n69), .B(n86), .C(n77), .D(n57), .E(n6319), .Z(
        n6318) );
  HS65_LL_NAND4ABX3 U15120 ( .A(n8370), .B(n8371), .C(n8372), .D(n8373), .Z(
        n2778) );
  HS65_LL_NAND4ABX3 U15121 ( .A(n8417), .B(n8418), .C(n8419), .D(n8420), .Z(
        n8370) );
  HS65_LL_OAI212X5 U15122 ( .A(n8415), .B(n7630), .C(n7677), .D(n7636), .E(
        n8416), .Z(n8371) );
  HS65_LL_AOI212X4 U15123 ( .A(n592), .B(n608), .C(n588), .D(n602), .E(n8374), 
        .Z(n8373) );
  HS65_LL_NAND4ABX3 U15124 ( .A(n4537), .B(n4538), .C(n4539), .D(n4540), .Z(
        n2771) );
  HS65_LL_NAND4ABX3 U15125 ( .A(n4573), .B(n4574), .C(n4575), .D(n4576), .Z(
        n4537) );
  HS65_LL_OAI212X5 U15126 ( .A(n4565), .B(n4566), .C(n4478), .D(n4567), .E(
        n4568), .Z(n4538) );
  HS65_LL_AOI212X4 U15127 ( .A(n9), .B(n34), .C(n30), .D(n14), .E(n4541), .Z(
        n4540) );
  HS65_LL_NAND4ABX3 U15128 ( .A(n6130), .B(n6131), .C(n6132), .D(n6133), .Z(
        n2763) );
  HS65_LL_NAND4ABX3 U15129 ( .A(n6166), .B(n6167), .C(n6168), .D(n6169), .Z(
        n6130) );
  HS65_LL_OAI212X5 U15130 ( .A(n6158), .B(n6159), .C(n6071), .D(n6160), .E(
        n6161), .Z(n6131) );
  HS65_LL_AOI212X4 U15131 ( .A(n531), .B(n556), .C(n552), .D(n536), .E(n6134), 
        .Z(n6133) );
  HS65_LL_OAI212X5 U15132 ( .A(n3808), .B(n2845), .C(n2995), .D(n3380), .E(
        n4041), .Z(n4039) );
  HS65_LL_CB4I1X9 U15133 ( .A(n3972), .B(n3204), .C(n3846), .D(n3809), .Z(
        n4041) );
  HS65_LL_NAND4ABX3 U15134 ( .A(n8156), .B(n8157), .C(n8158), .D(n8159), .Z(
        n2803) );
  HS65_LL_NAND4ABX3 U15135 ( .A(n8184), .B(n8185), .C(n8186), .D(n8187), .Z(
        n8156) );
  HS65_LL_OAI212X5 U15136 ( .A(n7658), .B(n8179), .C(n7869), .D(n7905), .E(
        n8180), .Z(n8157) );
  HS65_LL_NOR3AX2 U15137 ( .A(n8013), .B(n8162), .C(n8163), .Z(n8158) );
  HS65_LL_NAND4ABX3 U15138 ( .A(n8308), .B(n8309), .C(n8310), .D(n8311), .Z(
        n3002) );
  HS65_LL_NAND4ABX3 U15139 ( .A(n8365), .B(n8366), .C(n8367), .D(n8368), .Z(
        n8308) );
  HS65_LL_OAI212X5 U15140 ( .A(n8362), .B(n7943), .C(n7770), .D(n8363), .E(
        n8364), .Z(n8309) );
  HS65_LL_AOI212X4 U15141 ( .A(n323), .B(n339), .C(n329), .D(n344), .E(n8312), 
        .Z(n8311) );
  HS65_LL_NAND4ABX3 U15142 ( .A(n4761), .B(n4762), .C(n4763), .D(n4764), .Z(
        n2819) );
  HS65_LL_NAND4ABX3 U15143 ( .A(n4796), .B(n4797), .C(n4798), .D(n4799), .Z(
        n4761) );
  HS65_LL_OAI212X5 U15144 ( .A(n4788), .B(n4789), .C(n4493), .D(n4790), .E(
        n4791), .Z(n4762) );
  HS65_LL_AOI212X4 U15145 ( .A(n462), .B(n480), .C(n476), .D(n458), .E(n4765), 
        .Z(n4764) );
  HS65_LL_NAND4ABX3 U15146 ( .A(n6354), .B(n6355), .C(n6356), .D(n6357), .Z(
        n2811) );
  HS65_LL_NAND4ABX3 U15147 ( .A(n6389), .B(n6390), .C(n6391), .D(n6392), .Z(
        n6354) );
  HS65_LL_OAI212X5 U15148 ( .A(n6381), .B(n6382), .C(n6086), .D(n6383), .E(
        n6384), .Z(n6355) );
  HS65_LL_AOI212X4 U15149 ( .A(n287), .B(n305), .C(n301), .D(n283), .E(n6358), 
        .Z(n6357) );
  HS65_LL_NOR4ABX2 U15150 ( .A(n3902), .B(n3903), .C(n3904), .D(n3905), .Z(
        n2897) );
  HS65_LL_CBI4I1X5 U15151 ( .A(n3048), .B(n3251), .C(n2914), .D(n3624), .Z(
        n3904) );
  HS65_LL_AOI212X4 U15152 ( .A(n170), .B(n155), .C(n156), .D(n3912), .E(n3913), 
        .Z(n3902) );
  HS65_LL_CBI4I6X5 U15153 ( .A(n172), .B(n3597), .C(n157), .D(n3911), .Z(n3903) );
  HS65_LL_OAI212X5 U15154 ( .A(n3451), .B(n2940), .C(n2857), .D(n3096), .E(
        n3927), .Z(n3924) );
  HS65_LL_CB4I1X9 U15155 ( .A(n3928), .B(n2939), .C(n3491), .D(n3452), .Z(
        n3927) );
  HS65_LL_OAI212X5 U15156 ( .A(n5709), .B(n4485), .C(n5013), .D(n5026), .E(
        n5710), .Z(n5708) );
  HS65_LL_OAI21X3 U15157 ( .A(n24), .B(n17), .C(n40), .Z(n5710) );
  HS65_LL_NOR3X4 U15158 ( .A(n44), .B(n46), .C(n34), .Z(n5709) );
  HS65_LL_OAI212X5 U15159 ( .A(n7301), .B(n6078), .C(n6606), .D(n6619), .E(
        n7302), .Z(n7300) );
  HS65_LL_OAI21X3 U15160 ( .A(n546), .B(n539), .C(n562), .Z(n7302) );
  HS65_LL_NOR3X4 U15161 ( .A(n566), .B(n568), .C(n556), .Z(n7301) );
  HS65_LL_NAND4ABX3 U15162 ( .A(n3013), .B(n3014), .C(n3015), .D(n3016), .Z(
        n2638) );
  HS65_LL_NAND4ABX3 U15163 ( .A(n3049), .B(n3050), .C(n3051), .D(n3052), .Z(
        n3013) );
  HS65_LL_OAI212X5 U15164 ( .A(n3041), .B(n3042), .C(n3043), .D(n2918), .E(
        n3044), .Z(n3014) );
  HS65_LL_AOI212X4 U15165 ( .A(n142), .B(n167), .C(n147), .D(n164), .E(n3017), 
        .Z(n3016) );
  HS65_LL_OAI212X5 U15166 ( .A(n8832), .B(n7713), .C(n8473), .D(n8178), .E(
        n9091), .Z(n9089) );
  HS65_LL_CBI4I6X5 U15167 ( .A(n135), .B(n127), .C(n113), .D(n8829), .Z(n9091)
         );
  HS65_LL_OAI212X5 U15168 ( .A(n8742), .B(n7675), .C(n8421), .D(n8155), .E(
        n9033), .Z(n9031) );
  HS65_LL_CBI4I6X5 U15169 ( .A(n615), .B(n607), .C(n593), .D(n8739), .Z(n9033)
         );
  HS65_LL_NAND4ABX3 U15170 ( .A(n3164), .B(n3165), .C(n3166), .D(n3167), .Z(
        n2692) );
  HS65_LL_NAND4ABX3 U15171 ( .A(n3199), .B(n3200), .C(n3201), .D(n3202), .Z(
        n3164) );
  HS65_LL_OAI212X5 U15172 ( .A(n3191), .B(n3192), .C(n3193), .D(n2830), .E(
        n3194), .Z(n3165) );
  HS65_LL_AOI212X4 U15173 ( .A(n420), .B(n439), .C(n415), .D(n442), .E(n3168), 
        .Z(n3167) );
  HS65_LL_NAND4ABX3 U15174 ( .A(n3219), .B(n3220), .C(n3221), .D(n3222), .Z(
        n2645) );
  HS65_LL_OAI212X5 U15175 ( .A(n3278), .B(n3032), .C(n3279), .D(n3280), .E(
        n3281), .Z(n3220) );
  HS65_LL_NAND4ABX3 U15176 ( .A(n3282), .B(n3283), .C(n3284), .D(n3285), .Z(
        n3219) );
  HS65_LL_AOI212X4 U15177 ( .A(n156), .B(n171), .C(n180), .D(n151), .E(n3223), 
        .Z(n3222) );
  HS65_LL_NAND4ABX3 U15178 ( .A(n8845), .B(n8846), .C(n8847), .D(n8848), .Z(
        n3000) );
  HS65_LL_AOI212X4 U15179 ( .A(n324), .B(n350), .C(n323), .D(n8619), .E(n8870), 
        .Z(n8847) );
  HS65_LL_CBI4I1X5 U15180 ( .A(n8629), .B(n7769), .C(n7951), .D(n8872), .Z(
        n8846) );
  HS65_LL_CB4I6X9 U15181 ( .A(n355), .B(n349), .C(n330), .D(n8574), .Z(n8845)
         );
  HS65_LL_NOR4ABX2 U15182 ( .A(n3055), .B(n3056), .C(n3057), .D(n3058), .Z(
        n2651) );
  HS65_LL_NAND4ABX3 U15183 ( .A(n3063), .B(n3064), .C(n3065), .D(n3066), .Z(
        n3057) );
  HS65_LL_OAI212X5 U15184 ( .A(n3059), .B(n2956), .C(n3060), .D(n3061), .E(
        n3062), .Z(n3058) );
  HS65_LL_AOI212X4 U15185 ( .A(n201), .B(n208), .C(n226), .D(n196), .E(n3068), 
        .Z(n3056) );
  HS65_LL_NOR4ABX2 U15186 ( .A(n7955), .B(n7956), .C(n7957), .D(n7958), .Z(
        n2755) );
  HS65_LL_NAND4ABX3 U15187 ( .A(n7967), .B(n7968), .C(n7969), .D(n7970), .Z(
        n7957) );
  HS65_LL_OAI212X5 U15188 ( .A(n7959), .B(n7960), .C(n7961), .D(n7851), .E(
        n7962), .Z(n7958) );
  HS65_LL_AOI212X4 U15189 ( .A(n398), .B(n366), .C(n367), .D(n396), .E(n7972), 
        .Z(n7956) );
  HS65_LL_NAND4ABX3 U15190 ( .A(n2982), .B(n2983), .C(n2984), .D(n2985), .Z(
        n2687) );
  HS65_LL_CBI4I1X5 U15191 ( .A(n2993), .B(n2994), .C(n2995), .D(n2996), .Z(
        n2983) );
  HS65_LL_AOI212X4 U15192 ( .A(n417), .B(n433), .C(n412), .D(n428), .E(n2991), 
        .Z(n2984) );
  HS65_LL_CBI4I1X5 U15193 ( .A(n2997), .B(n2830), .C(n2998), .D(n2999), .Z(
        n2982) );
  HS65_LL_IVX9 U15194 ( .A(n8005), .Z(n615) );
  HS65_LL_OAI212X5 U15195 ( .A(n8081), .B(n8082), .C(n7960), .D(n8067), .E(
        n8083), .Z(n8070) );
  HS65_LL_OAI21X3 U15196 ( .A(n372), .B(n366), .C(n400), .Z(n8083) );
  HS65_LL_NOR2X6 U15197 ( .A(n375), .B(n377), .Z(n8081) );
  HS65_LL_OAI212X5 U15198 ( .A(n3449), .B(n3450), .C(n3451), .D(n3114), .E(
        n3452), .Z(n3438) );
  HS65_LL_NOR2X6 U15199 ( .A(n199), .B(n202), .Z(n3449) );
  HS65_LL_OAI212X5 U15200 ( .A(n3032), .B(n3033), .C(n3034), .D(n3035), .E(
        n3036), .Z(n3022) );
  HS65_LL_OAI21X3 U15201 ( .A(n158), .B(n157), .C(n172), .Z(n3036) );
  HS65_LL_NOR4ABX2 U15202 ( .A(n8124), .B(n8125), .C(n8126), .D(n8127), .Z(
        n2779) );
  HS65_LL_NAND4ABX3 U15203 ( .A(n8133), .B(n8134), .C(n8135), .D(n8136), .Z(
        n8126) );
  HS65_LL_OAI212X5 U15204 ( .A(n7637), .B(n8128), .C(n7806), .D(n7807), .E(
        n8129), .Z(n8127) );
  HS65_LL_NOR3AX2 U15205 ( .A(n8000), .B(n8139), .C(n8140), .Z(n8124) );
  HS65_LL_IVX9 U15206 ( .A(n4093), .Z(n163) );
  HS65_LL_NOR4ABX2 U15207 ( .A(n4722), .B(n4723), .C(n4724), .D(n4725), .Z(
        n2795) );
  HS65_LL_NAND4ABX3 U15208 ( .A(n4735), .B(n4736), .C(n4737), .D(n4738), .Z(
        n4724) );
  HS65_LL_OAI212X5 U15209 ( .A(n4726), .B(n4727), .C(n4454), .D(n4728), .E(
        n4729), .Z(n4725) );
  HS65_LL_AOI212X4 U15210 ( .A(n245), .B(n263), .C(n259), .D(n241), .E(n4739), 
        .Z(n4723) );
  HS65_LL_NAND4ABX3 U15211 ( .A(n6397), .B(n6398), .C(n6399), .D(n6400), .Z(
        n3205) );
  HS65_LL_NAND4ABX3 U15212 ( .A(n6457), .B(n6458), .C(n6459), .D(n6460), .Z(
        n6397) );
  HS65_LL_OAI212X5 U15213 ( .A(n6453), .B(n6219), .C(n6454), .D(n6455), .E(
        n6456), .Z(n6398) );
  HS65_LL_AOI212X4 U15214 ( .A(n498), .B(n517), .C(n526), .D(n501), .E(n6401), 
        .Z(n6400) );
  HS65_LL_NAND4ABX3 U15215 ( .A(n4804), .B(n4805), .C(n4806), .D(n4807), .Z(
        n3213) );
  HS65_LL_NAND4ABX3 U15216 ( .A(n4864), .B(n4865), .C(n4866), .D(n4867), .Z(
        n4804) );
  HS65_LL_OAI212X5 U15217 ( .A(n4860), .B(n4626), .C(n4861), .D(n4862), .E(
        n4863), .Z(n4805) );
  HS65_LL_AOI212X4 U15218 ( .A(n674), .B(n693), .C(n702), .D(n677), .E(n4808), 
        .Z(n4807) );
  HS65_LL_IVX9 U15219 ( .A(n3270), .Z(n147) );
  HS65_LL_OAI212X5 U15220 ( .A(n4116), .B(n3053), .C(n3588), .D(n3269), .E(
        n4117), .Z(n4115) );
  HS65_LL_NOR3X4 U15221 ( .A(n167), .B(n177), .C(n179), .Z(n4116) );
  HS65_LL_OAI21X3 U15222 ( .A(n153), .B(n149), .C(n173), .Z(n4117) );
  HS65_LL_OAI212X5 U15223 ( .A(n8526), .B(n8527), .C(n8528), .D(n7768), .E(
        n8529), .Z(n8515) );
  HS65_LL_NOR2X6 U15224 ( .A(n328), .B(n325), .Z(n8526) );
  HS65_LL_OAI212X5 U15225 ( .A(n3573), .B(n3574), .C(n3575), .D(n3270), .E(
        n3576), .Z(n3562) );
  HS65_LL_NOR2X6 U15226 ( .A(n154), .B(n157), .Z(n3573) );
  HS65_LL_NOR4ABX2 U15227 ( .A(n3978), .B(n3979), .C(n3980), .D(n3981), .Z(
        n2896) );
  HS65_LL_CBI4I1X5 U15228 ( .A(n3048), .B(n3984), .C(n3035), .D(n3633), .Z(
        n3980) );
  HS65_LL_CBI4I1X5 U15229 ( .A(n2919), .B(n3982), .C(n3270), .D(n3983), .Z(
        n3981) );
  HS65_LL_AOI222X2 U15230 ( .A(n148), .B(n167), .C(n156), .D(n3995), .E(n152), 
        .F(n163), .Z(n3978) );
  HS65_LL_OAI212X5 U15231 ( .A(n7820), .B(n7632), .C(n7821), .D(n7822), .E(
        n7823), .Z(n7819) );
  HS65_LL_NOR3X4 U15232 ( .A(n599), .B(n604), .C(n603), .Z(n7820) );
  HS65_LL_OAI21X3 U15233 ( .A(n585), .B(n580), .C(n611), .Z(n7823) );
  HS65_LL_OAI212X5 U15234 ( .A(n5622), .B(n4499), .C(n4610), .D(n5380), .E(
        n5623), .Z(n5621) );
  HS65_LL_NOR3X4 U15235 ( .A(n480), .B(n467), .C(n472), .Z(n5622) );
  HS65_LL_OAI21X3 U15236 ( .A(n451), .B(n460), .C(n482), .Z(n5623) );
  HS65_LL_OAI212X5 U15237 ( .A(n5597), .B(n4460), .C(n4593), .D(n5265), .E(
        n5598), .Z(n5596) );
  HS65_LL_NOR3X4 U15238 ( .A(n263), .B(n250), .C(n255), .Z(n5597) );
  HS65_LL_OAI21X3 U15239 ( .A(n234), .B(n243), .C(n265), .Z(n5598) );
  HS65_LL_OAI212X5 U15240 ( .A(n7214), .B(n6092), .C(n6203), .D(n6972), .E(
        n7215), .Z(n7213) );
  HS65_LL_NOR3X4 U15241 ( .A(n305), .B(n292), .C(n297), .Z(n7214) );
  HS65_LL_OAI21X3 U15242 ( .A(n276), .B(n285), .C(n307), .Z(n7215) );
  HS65_LL_OAI212X5 U15243 ( .A(n5771), .B(n4525), .C(n5135), .D(n5148), .E(
        n5772), .Z(n5770) );
  HS65_LL_NOR3X4 U15244 ( .A(n689), .B(n701), .C(n699), .Z(n5771) );
  HS65_LL_OAI21X3 U15245 ( .A(n679), .B(n672), .C(n695), .Z(n5772) );
  HS65_LL_OAI212X5 U15246 ( .A(n7363), .B(n6118), .C(n6727), .D(n6740), .E(
        n7364), .Z(n7362) );
  HS65_LL_NOR3X4 U15247 ( .A(n513), .B(n525), .C(n523), .Z(n7363) );
  HS65_LL_OAI21X3 U15248 ( .A(n503), .B(n496), .C(n519), .Z(n7364) );
  HS65_LL_IVX9 U15249 ( .A(n2917), .Z(n157) );
  HS65_LL_NAND4ABX3 U15250 ( .A(n5483), .B(n5484), .C(n5485), .D(n5486), .Z(
        n3211) );
  HS65_LL_CBI4I1X5 U15251 ( .A(n4649), .B(n4848), .C(n4847), .D(n5168), .Z(
        n5483) );
  HS65_LL_AOI212X4 U15252 ( .A(n673), .B(n692), .C(n674), .D(n5492), .E(n5493), 
        .Z(n5485) );
  HS65_LL_CBI4I1X5 U15253 ( .A(n5494), .B(n4850), .C(n4533), .D(n5495), .Z(
        n5484) );
  HS65_LL_NAND4ABX3 U15254 ( .A(n7075), .B(n7076), .C(n7077), .D(n7078), .Z(
        n3008) );
  HS65_LL_CBI4I1X5 U15255 ( .A(n6242), .B(n6441), .C(n6440), .D(n6760), .Z(
        n7075) );
  HS65_LL_AOI212X4 U15256 ( .A(n497), .B(n516), .C(n498), .D(n7084), .E(n7085), 
        .Z(n7077) );
  HS65_LL_CBI4I1X5 U15257 ( .A(n7086), .B(n6443), .C(n6126), .D(n7087), .Z(
        n7076) );
  HS65_LL_IVX9 U15258 ( .A(n3033), .Z(n170) );
  HS65_LL_NAND2X7 U15259 ( .A(n7965), .B(n7859), .Z(n8080) );
  HS65_LL_NOR2X6 U15260 ( .A(n3054), .B(n3035), .Z(n3654) );
  HS65_LL_IVX9 U15261 ( .A(n6727), .Z(n498) );
  HS65_LL_IVX9 U15262 ( .A(n5135), .Z(n674) );
  HS65_LL_IVX9 U15263 ( .A(n5148), .Z(n691) );
  HS65_LL_NAND2X7 U15264 ( .A(n8033), .B(n7941), .Z(n8324) );
  HS65_LL_IVX9 U15265 ( .A(n3574), .Z(n175) );
  HS65_LL_OAI212X5 U15266 ( .A(n6277), .B(n6278), .C(n6076), .D(n6159), .E(
        n6279), .Z(n6266) );
  HS65_LL_NOR2X6 U15267 ( .A(n545), .B(n544), .Z(n6277) );
  HS65_LL_OAI21X3 U15268 ( .A(n542), .B(n531), .C(n557), .Z(n6279) );
  HS65_LL_OAI212X5 U15269 ( .A(n4684), .B(n4685), .C(n4483), .D(n4566), .E(
        n4686), .Z(n4673) );
  HS65_LL_NOR2X6 U15270 ( .A(n23), .B(n22), .Z(n4684) );
  HS65_LL_OAI21X3 U15271 ( .A(n20), .B(n9), .C(n35), .Z(n4686) );
  HS65_LL_AOI212X4 U15272 ( .A(n16), .B(n28), .C(n41), .D(n25), .E(n5716), .Z(
        n5715) );
  HS65_LL_CBI4I1X5 U15273 ( .A(n4552), .B(n4478), .C(n4567), .D(n5110), .Z(
        n5716) );
  HS65_LL_AOI212X4 U15274 ( .A(n538), .B(n550), .C(n563), .D(n547), .E(n7308), 
        .Z(n7307) );
  HS65_LL_CBI4I1X5 U15275 ( .A(n6145), .B(n6071), .C(n6160), .D(n6703), .Z(
        n7308) );
  HS65_LL_NOR2X6 U15276 ( .A(n3982), .B(n2917), .Z(n3611) );
  HS65_LL_NOR2X6 U15277 ( .A(n3253), .B(n3035), .Z(n3655) );
  HS65_LL_NOR2X6 U15278 ( .A(n7980), .B(n7850), .Z(n8217) );
  HS65_LL_IVX9 U15279 ( .A(n5572), .Z(n697) );
  HS65_LL_AOI212X4 U15280 ( .A(n242), .B(n254), .C(n267), .D(n235), .E(n5834), 
        .Z(n5832) );
  HS65_LL_CBI4I1X5 U15281 ( .A(n4733), .B(n4454), .C(n4728), .D(n5331), .Z(
        n5834) );
  HS65_LL_AOI212X4 U15282 ( .A(n459), .B(n471), .C(n484), .D(n452), .E(n5893), 
        .Z(n5891) );
  HS65_LL_CBI4I1X5 U15283 ( .A(n4775), .B(n4493), .C(n4790), .D(n5446), .Z(
        n5893) );
  HS65_LL_AOI212X4 U15284 ( .A(n671), .B(n683), .C(n696), .D(n680), .E(n5778), 
        .Z(n5776) );
  HS65_LL_CBI4I1X5 U15285 ( .A(n4629), .B(n4534), .C(n4644), .D(n5215), .Z(
        n5778) );
  HS65_LL_AOI212X4 U15286 ( .A(n284), .B(n296), .C(n309), .D(n277), .E(n7485), 
        .Z(n7483) );
  HS65_LL_CBI4I1X5 U15287 ( .A(n6368), .B(n6086), .C(n6383), .D(n7038), .Z(
        n7485) );
  HS65_LL_AOI212X4 U15288 ( .A(n495), .B(n507), .C(n520), .D(n504), .E(n7370), 
        .Z(n7368) );
  HS65_LL_CBI4I1X5 U15289 ( .A(n6222), .B(n6127), .C(n6237), .D(n6807), .Z(
        n7370) );
  HS65_LL_AOI212X4 U15290 ( .A(n54), .B(n72), .C(n81), .D(n66), .E(n7426), .Z(
        n7424) );
  HS65_LL_CBI4I1X5 U15291 ( .A(n6329), .B(n6047), .C(n6344), .D(n6923), .Z(
        n7426) );
  HS65_LL_NOR2X6 U15292 ( .A(n7846), .B(n7751), .Z(n8265) );
  HS65_LL_NOR2X6 U15293 ( .A(n5555), .B(n5630), .Z(n5460) );
  HS65_LL_NOR2X6 U15294 ( .A(n5571), .B(n5581), .Z(n5230) );
  HS65_LL_NOR2X6 U15295 ( .A(n7163), .B(n7173), .Z(n6822) );
  HS65_LL_NOR2X6 U15296 ( .A(n8630), .B(n8033), .Z(n8566) );
  HS65_LL_NOR2X6 U15297 ( .A(n8155), .B(n7636), .Z(n8384) );
  HS65_LL_OAI212X5 U15298 ( .A(n8413), .B(n7783), .C(n7836), .D(n8128), .E(
        n8414), .Z(n8404) );
  HS65_LL_NOR2X6 U15299 ( .A(n586), .B(n588), .Z(n8413) );
  HS65_LL_OAI21X3 U15300 ( .A(n593), .B(n584), .C(n607), .Z(n8414) );
  HS65_LL_OAI212X5 U15301 ( .A(n8465), .B(n7882), .C(n7875), .D(n8179), .E(
        n8466), .Z(n8456) );
  HS65_LL_NOR2X6 U15302 ( .A(n106), .B(n108), .Z(n8465) );
  HS65_LL_OAI21X3 U15303 ( .A(n113), .B(n104), .C(n127), .Z(n8466) );
  HS65_LL_IVX9 U15304 ( .A(n7170), .Z(n510) );
  HS65_LL_IVX9 U15305 ( .A(n5578), .Z(n686) );
  HS65_LL_NAND2X7 U15306 ( .A(n8132), .B(n7835), .Z(n8385) );
  HS65_LL_NAND2X7 U15307 ( .A(n8183), .B(n7874), .Z(n8437) );
  HS65_LL_NOR2X6 U15308 ( .A(n3069), .B(n3464), .Z(n3505) );
  HS65_LL_NOR2X6 U15309 ( .A(n2838), .B(n2992), .Z(n3859) );
  HS65_LL_AOI212X4 U15310 ( .A(n96), .B(n118), .C(n107), .D(n130), .E(n7904), 
        .Z(n7903) );
  HS65_LL_CBI4I1X5 U15311 ( .A(n7664), .B(n7869), .C(n7905), .D(n7906), .Z(
        n7904) );
  HS65_LL_AOI212X4 U15312 ( .A(n576), .B(n598), .C(n587), .D(n610), .E(n7805), 
        .Z(n7804) );
  HS65_LL_CBI4I1X5 U15313 ( .A(n7624), .B(n7806), .C(n7807), .D(n7808), .Z(
        n7805) );
  HS65_LL_NOR2X6 U15314 ( .A(n6236), .B(n7164), .Z(n6434) );
  HS65_LL_NOR2X6 U15315 ( .A(n4643), .B(n5572), .Z(n4841) );
  HS65_LL_NOR2X6 U15316 ( .A(n7099), .B(n7094), .Z(n6687) );
  HS65_LL_NOR2X6 U15317 ( .A(n5507), .B(n5502), .Z(n5094) );
  HS65_LL_IVX9 U15318 ( .A(n3032), .Z(n143) );
  HS65_LL_NOR2X6 U15319 ( .A(n8048), .B(n7951), .Z(n8606) );
  HS65_LL_NAND2X7 U15320 ( .A(n4732), .B(n4461), .Z(n4897) );
  HS65_LL_NAND2X7 U15321 ( .A(n4794), .B(n4500), .Z(n4950) );
  HS65_LL_NAND2X7 U15322 ( .A(n6387), .B(n6093), .Z(n6543) );
  HS65_LL_NAND2X7 U15323 ( .A(n6348), .B(n6054), .Z(n6490) );
  HS65_LL_NAND2X7 U15324 ( .A(n6241), .B(n7088), .Z(n6415) );
  HS65_LL_NAND2X7 U15325 ( .A(n4648), .B(n5496), .Z(n4822) );
  HS65_LL_NOR2X6 U15326 ( .A(n4789), .B(n5380), .Z(n5457) );
  HS65_LL_NOR2X6 U15327 ( .A(n4643), .B(n5148), .Z(n5227) );
  HS65_LL_NOR2X6 U15328 ( .A(n6236), .B(n6740), .Z(n6819) );
  HS65_LL_NOR2X6 U15329 ( .A(n4493), .B(n5629), .Z(n4782) );
  HS65_LL_NOR2X6 U15330 ( .A(n4454), .B(n5604), .Z(n4755) );
  HS65_LL_NOR2X6 U15331 ( .A(n6086), .B(n7221), .Z(n6375) );
  HS65_LL_NOR2X6 U15332 ( .A(n4534), .B(n5578), .Z(n4636) );
  HS65_LL_NOR2X6 U15333 ( .A(n6127), .B(n7170), .Z(n6229) );
  HS65_LL_NOR2X6 U15334 ( .A(n6047), .B(n7196), .Z(n6336) );
  HS65_LL_NOR2X6 U15335 ( .A(n6164), .B(n6261), .Z(n6656) );
  HS65_LL_NOR2X6 U15336 ( .A(n4571), .B(n4668), .Z(n5063) );
  HS65_LL_NOR2X6 U15337 ( .A(n4478), .B(n5514), .Z(n4559) );
  HS65_LL_NOR2X6 U15338 ( .A(n6071), .B(n7106), .Z(n6152) );
  HS65_LL_NOR2X6 U15339 ( .A(n3807), .B(n3192), .Z(n3378) );
  HS65_LL_NOR2X6 U15340 ( .A(n2913), .B(n3253), .Z(n3627) );
  HS65_LL_NOR2X6 U15341 ( .A(n8128), .B(n7633), .Z(n7799) );
  HS65_LL_NOR2X6 U15342 ( .A(n8179), .B(n7653), .Z(n7898) );
  HS65_LL_NOR2X6 U15343 ( .A(n4566), .B(n5508), .Z(n4703) );
  HS65_LL_NOR2X6 U15344 ( .A(n6159), .B(n7100), .Z(n6296) );
  HS65_LL_NOR2X6 U15345 ( .A(n3692), .B(n3128), .Z(n3324) );
  HS65_LL_OAI212X5 U15346 ( .A(n3806), .B(n3807), .C(n3808), .D(n3396), .E(
        n3809), .Z(n3796) );
  HS65_LL_NOR2X6 U15347 ( .A(n412), .B(n408), .Z(n3806) );
  HS65_LL_NOR2X6 U15348 ( .A(n2913), .B(n3054), .Z(n3274) );
  HS65_LL_NOR2X6 U15349 ( .A(n2913), .B(n4093), .Z(n3608) );
  HS65_LL_OAI212X5 U15350 ( .A(n8554), .B(n8058), .C(n7949), .D(n7952), .E(
        n8555), .Z(n8544) );
  HS65_LL_NOR2X6 U15351 ( .A(n335), .B(n8498), .Z(n8554) );
  HS65_LL_OAI212X5 U15352 ( .A(n6618), .B(n6619), .C(n6261), .D(n6071), .E(
        n6620), .Z(n6608) );
  HS65_LL_NOR2X6 U15353 ( .A(n538), .B(n6593), .Z(n6618) );
  HS65_LL_OAI212X5 U15354 ( .A(n5025), .B(n5026), .C(n4668), .D(n4478), .E(
        n5027), .Z(n5015) );
  HS65_LL_NOR2X6 U15355 ( .A(n16), .B(n5000), .Z(n5025) );
  HS65_LL_NOR2X6 U15356 ( .A(n8028), .B(n8339), .Z(n8593) );
  HS65_LL_NOR2X6 U15357 ( .A(n7652), .B(n7662), .Z(n7924) );
  HS65_LL_NOR2X6 U15358 ( .A(n7632), .B(n7622), .Z(n7826) );
  HS65_LL_OAI212X5 U15359 ( .A(n3613), .B(n3269), .C(n2915), .D(n2918), .E(
        n3614), .Z(n3603) );
  HS65_LL_NOR2X6 U15360 ( .A(n150), .B(n3541), .Z(n3613) );
  HS65_LL_NOR2X6 U15361 ( .A(n8183), .B(n8473), .Z(n7728) );
  HS65_LL_NOR2X6 U15362 ( .A(n7951), .B(n7942), .Z(n8549) );
  HS65_LL_NOR2X6 U15363 ( .A(n3450), .B(n2926), .Z(n3094) );
  HS65_LL_NOR2X6 U15364 ( .A(n8178), .B(n8018), .Z(n8448) );
  HS65_LL_NOR2X6 U15365 ( .A(n8155), .B(n8005), .Z(n8396) );
  HS65_LL_NOR2X6 U15366 ( .A(n7992), .B(n7993), .Z(n7747) );
  HS65_LL_NOR2X6 U15367 ( .A(n3225), .B(n4093), .Z(n3246) );
  HS65_LL_NOR2X6 U15368 ( .A(n7846), .B(n8067), .Z(n8111) );
  HS65_LL_NAND2X7 U15369 ( .A(n3450), .B(n2857), .Z(n3101) );
  HS65_LL_NAND2X7 U15370 ( .A(n3043), .B(n4093), .Z(n3597) );
  HS65_LL_NOR2X6 U15371 ( .A(n3112), .B(n2932), .Z(n3523) );
  HS65_LL_NAND2X7 U15372 ( .A(n6164), .B(n7064), .Z(n6276) );
  HS65_LL_NAND2X7 U15373 ( .A(n4571), .B(n5472), .Z(n4683) );
  HS65_LL_NOR2X6 U15374 ( .A(n4485), .B(n5501), .Z(n5043) );
  HS65_LL_NOR2X6 U15375 ( .A(n6078), .B(n7093), .Z(n6636) );
  HS65_LL_NOR2X6 U15376 ( .A(n4661), .B(n4711), .Z(n4693) );
  HS65_LL_NOR2X6 U15377 ( .A(n6254), .B(n6304), .Z(n6286) );
  HS65_LL_NOR2X6 U15378 ( .A(n2855), .B(n2958), .Z(n2951) );
  HS65_LL_NAND2X7 U15379 ( .A(n8302), .B(n7848), .Z(n8110) );
  HS65_LL_NOR2X6 U15380 ( .A(n7664), .B(n7882), .Z(n8804) );
  HS65_LL_NOR2X6 U15381 ( .A(n7624), .B(n7783), .Z(n8714) );
  HS65_LL_NOR2X6 U15382 ( .A(n8397), .B(n7783), .Z(n8725) );
  HS65_LL_NAND2X7 U15383 ( .A(n5616), .B(n4995), .Z(n4980) );
  HS65_LL_NAND2X7 U15384 ( .A(n5572), .B(n4869), .Z(n4854) );
  HS65_LL_NAND2X7 U15385 ( .A(n7208), .B(n6588), .Z(n6573) );
  HS65_LL_NAND2X7 U15386 ( .A(n7164), .B(n6462), .Z(n6447) );
  HS65_LL_NOR2X6 U15387 ( .A(n7920), .B(n8179), .Z(n8816) );
  HS65_LL_NOR2X6 U15388 ( .A(n7822), .B(n8128), .Z(n8726) );
  HS65_LL_NOR2X6 U15389 ( .A(n7088), .B(n7171), .Z(n6753) );
  HS65_LL_NOR2X6 U15390 ( .A(n5496), .B(n5579), .Z(n5161) );
  HS65_LL_NOR2X6 U15391 ( .A(n4727), .B(n5533), .Z(n4907) );
  HS65_LL_NOR2X6 U15392 ( .A(n6343), .B(n7125), .Z(n6500) );
  HS65_LL_NOR2X6 U15393 ( .A(n6236), .B(n7163), .Z(n6425) );
  HS65_LL_NOR2X6 U15394 ( .A(n4643), .B(n5571), .Z(n4832) );
  HS65_LL_NOR2X6 U15395 ( .A(n8057), .B(n8058), .Z(n7765) );
  HS65_LL_NOR2X6 U15396 ( .A(n4876), .B(n4923), .Z(n4906) );
  HS65_LL_NOR2X6 U15397 ( .A(n4988), .B(n4976), .Z(n4959) );
  HS65_LL_NOR2X6 U15398 ( .A(n6581), .B(n6569), .Z(n6552) );
  HS65_LL_NOR2X6 U15399 ( .A(n6469), .B(n6516), .Z(n6499) );
  HS65_LL_NOR2X6 U15400 ( .A(n6455), .B(n6442), .Z(n6424) );
  HS65_LL_NOR2X6 U15401 ( .A(n4862), .B(n4849), .Z(n4831) );
  HS65_LL_NOR2X6 U15402 ( .A(n2932), .B(n2938), .Z(n3526) );
  HS65_LL_NOR2X6 U15403 ( .A(n2993), .B(n3185), .Z(n3178) );
  HS65_LL_NOR2X6 U15404 ( .A(n2968), .B(n3158), .Z(n3152) );
  HS65_LL_NOR2X6 U15405 ( .A(n3286), .B(n3994), .Z(n3566) );
  HS65_LL_NOR2X6 U15406 ( .A(n2913), .B(n3048), .Z(n3245) );
  HS65_LL_NOR2X6 U15407 ( .A(n3053), .B(n3048), .Z(n3630) );
  HS65_LL_IVX9 U15408 ( .A(n3043), .Z(n177) );
  HS65_LL_NOR2X6 U15409 ( .A(n7947), .B(n7940), .Z(n8337) );
  HS65_LL_NOR2X6 U15410 ( .A(n2272), .B(n2308), .Z(n2316) );
  HS65_LL_NOR2X6 U15411 ( .A(n1520), .B(n1556), .Z(n1564) );
  HS65_LL_NOR2X6 U15412 ( .A(n1896), .B(n1932), .Z(n1940) );
  HS65_LL_NOR2X6 U15413 ( .A(n5604), .B(n4882), .Z(n5306) );
  HS65_LL_NOR2X6 U15414 ( .A(n5629), .B(n4994), .Z(n5421) );
  HS65_LL_NOR2X6 U15415 ( .A(n5578), .B(n4868), .Z(n5190) );
  HS65_LL_NOR2X6 U15416 ( .A(n7221), .B(n6587), .Z(n7013) );
  HS65_LL_NOR2X6 U15417 ( .A(n7170), .B(n6461), .Z(n6782) );
  HS65_LL_NOR2X6 U15418 ( .A(n3970), .B(n3197), .Z(n3857) );
  HS65_LL_NOR2X6 U15419 ( .A(n3926), .B(n2931), .Z(n3502) );
  HS65_LL_NOR2X6 U15420 ( .A(n6142), .B(n7064), .Z(n6632) );
  HS65_LL_NOR2X6 U15421 ( .A(n4549), .B(n5472), .Z(n5039) );
  HS65_LL_NOR2X6 U15422 ( .A(n4549), .B(n4477), .Z(n5098) );
  HS65_LL_NOR2X6 U15423 ( .A(n6142), .B(n6070), .Z(n6691) );
  HS65_LL_NOR2X6 U15424 ( .A(n3095), .B(n2926), .Z(n3530) );
  HS65_LL_NOR2X6 U15425 ( .A(n4500), .B(n4773), .Z(n5394) );
  HS65_LL_NOR2X6 U15426 ( .A(n6093), .B(n6366), .Z(n6986) );
  HS65_LL_NOR2X6 U15427 ( .A(n5496), .B(n4627), .Z(n5162) );
  HS65_LL_NOR2X6 U15428 ( .A(n7088), .B(n6220), .Z(n6754) );
  HS65_LL_NOR2X6 U15429 ( .A(n3053), .B(n3982), .Z(n3626) );
  HS65_LL_NOR2X6 U15430 ( .A(n6303), .B(n7099), .Z(n6660) );
  HS65_LL_NOR2X6 U15431 ( .A(n4710), .B(n5507), .Z(n5067) );
  HS65_LL_NOR2X6 U15432 ( .A(n6440), .B(n7163), .Z(n6781) );
  HS65_LL_NOR2X6 U15433 ( .A(n4847), .B(n5571), .Z(n5189) );
  HS65_LL_NOR2X6 U15434 ( .A(n4975), .B(n5555), .Z(n5420) );
  HS65_LL_NOR2X6 U15435 ( .A(n4922), .B(n5533), .Z(n5305) );
  HS65_LL_NOR2X6 U15436 ( .A(n6568), .B(n7147), .Z(n7012) );
  HS65_LL_NOR2X6 U15437 ( .A(n6515), .B(n7125), .Z(n6897) );
  HS65_LL_AOI212X4 U15438 ( .A(n241), .B(n251), .C(n264), .D(n5333), .E(n4464), 
        .Z(n5323) );
  HS65_LL_NAND2X7 U15439 ( .A(n4586), .B(n4923), .Z(n5333) );
  HS65_LL_IVX9 U15440 ( .A(n5334), .Z(n251) );
  HS65_LL_AOI212X4 U15441 ( .A(n458), .B(n468), .C(n481), .D(n5448), .E(n4503), 
        .Z(n5438) );
  HS65_LL_NAND2X7 U15442 ( .A(n4603), .B(n4976), .Z(n5448) );
  HS65_LL_IVX9 U15443 ( .A(n5449), .Z(n468) );
  HS65_LL_AOI212X4 U15444 ( .A(n669), .B(n687), .C(n697), .D(n5217), .E(n5218), 
        .Z(n5207) );
  HS65_LL_NAND2X7 U15445 ( .A(n4533), .B(n4849), .Z(n5217) );
  HS65_LL_IVX9 U15446 ( .A(n5219), .Z(n687) );
  HS65_LL_AOI212X4 U15447 ( .A(n283), .B(n293), .C(n306), .D(n7040), .E(n6096), 
        .Z(n7030) );
  HS65_LL_NAND2X7 U15448 ( .A(n6196), .B(n6569), .Z(n7040) );
  HS65_LL_IVX9 U15449 ( .A(n7041), .Z(n293) );
  HS65_LL_AOI212X4 U15450 ( .A(n493), .B(n511), .C(n521), .D(n6809), .E(n6810), 
        .Z(n6799) );
  HS65_LL_NAND2X7 U15451 ( .A(n6126), .B(n6442), .Z(n6809) );
  HS65_LL_IVX9 U15452 ( .A(n6811), .Z(n511) );
  HS65_LL_AOI212X4 U15453 ( .A(n99), .B(n121), .C(n132), .D(n8831), .E(n7877), 
        .Z(n8823) );
  HS65_LL_NAND2X7 U15454 ( .A(n7724), .B(n8178), .Z(n8831) );
  HS65_LL_IVX9 U15455 ( .A(n8832), .Z(n121) );
  HS65_LL_NOR2X6 U15456 ( .A(n5616), .B(n5630), .Z(n5434) );
  HS65_LL_NOR2X6 U15457 ( .A(n5572), .B(n5581), .Z(n5203) );
  HS65_LL_NOR2X6 U15458 ( .A(n7164), .B(n7173), .Z(n6795) );
  HS65_LL_NOR2X6 U15459 ( .A(n7870), .B(n7724), .Z(n8788) );
  HS65_LL_NOR2X6 U15460 ( .A(n7831), .B(n7686), .Z(n8698) );
  HS65_LL_NOR2X6 U15461 ( .A(n8369), .B(n8048), .Z(n8552) );
  HS65_LL_NOR2X6 U15462 ( .A(n6145), .B(n6254), .Z(n6663) );
  HS65_LL_NOR2X6 U15463 ( .A(n4552), .B(n4661), .Z(n5070) );
  HS65_LL_NAND2X7 U15464 ( .A(n5508), .B(n4668), .Z(n4716) );
  HS65_LL_NAND2X7 U15465 ( .A(n7653), .B(n8473), .Z(n7928) );
  HS65_LL_NAND2X7 U15466 ( .A(n7633), .B(n8421), .Z(n7830) );
  HS65_LL_NAND2X7 U15467 ( .A(n7100), .B(n6261), .Z(n6309) );
  HS65_LL_NOR2X6 U15468 ( .A(n3615), .B(n3574), .Z(n3587) );
  HS65_LL_NOR2X6 U15469 ( .A(n8313), .B(n7943), .Z(n8344) );
  HS65_LL_NAND2X7 U15470 ( .A(n8527), .B(n7949), .Z(n8343) );
  HS65_LL_NOR2X6 U15471 ( .A(n7846), .B(n7858), .Z(n8104) );
  HS65_LL_NOR2X6 U15472 ( .A(n3252), .B(n3280), .Z(n3234) );
  HS65_LL_NAND2X7 U15473 ( .A(n3574), .B(n2915), .Z(n3257) );
  HS65_LL_NOR2X6 U15474 ( .A(n4670), .B(n4484), .Z(n4704) );
  HS65_LL_NOR2X6 U15475 ( .A(n6263), .B(n6077), .Z(n6297) );
  HS65_LL_NAND2X7 U15476 ( .A(n7630), .B(n8397), .Z(n8130) );
  HS65_LL_NAND2X7 U15477 ( .A(n7650), .B(n8449), .Z(n8181) );
  HS65_LL_NOR2X6 U15478 ( .A(n4552), .B(n5501), .Z(n5060) );
  HS65_LL_NOR2X6 U15479 ( .A(n6145), .B(n7093), .Z(n6653) );
  HS65_LL_NOR2X6 U15480 ( .A(n2830), .B(n3406), .Z(n3779) );
  HS65_LL_NOR2X6 U15481 ( .A(n4794), .B(n4995), .Z(n5416) );
  HS65_LL_NOR2X6 U15482 ( .A(n6387), .B(n6588), .Z(n7008) );
  HS65_LL_NOR2X6 U15483 ( .A(n4732), .B(n4883), .Z(n5301) );
  HS65_LL_NOR2X6 U15484 ( .A(n4648), .B(n4869), .Z(n5185) );
  HS65_LL_NOR2X6 U15485 ( .A(n6241), .B(n6462), .Z(n6777) );
  HS65_LL_NOR2X6 U15486 ( .A(n3095), .B(n2931), .Z(n3429) );
  HS65_LL_NOR2X6 U15487 ( .A(n8123), .B(n7980), .Z(n8251) );
  HS65_LL_NOR2X6 U15488 ( .A(n3271), .B(n3982), .Z(n3631) );
  HS65_LL_NOR2X6 U15489 ( .A(n4566), .B(n5507), .Z(n4694) );
  HS65_LL_NOR2X6 U15490 ( .A(n6159), .B(n7099), .Z(n6287) );
  HS65_LL_NOR2X6 U15491 ( .A(n7835), .B(n7619), .Z(n7798) );
  HS65_LL_NOR2X6 U15492 ( .A(n7874), .B(n7656), .Z(n7897) );
  HS65_LL_NOR2X6 U15493 ( .A(n7064), .B(n7093), .Z(n6633) );
  HS65_LL_NOR2X6 U15494 ( .A(n5472), .B(n5501), .Z(n5040) );
  HS65_LL_NOR2X6 U15495 ( .A(n8369), .B(n8630), .Z(n8594) );
  HS65_LL_NOR2X6 U15496 ( .A(n8005), .B(n7675), .Z(n8393) );
  HS65_LL_NOR2X6 U15497 ( .A(n8018), .B(n7713), .Z(n8445) );
  HS65_LL_NOR2X6 U15498 ( .A(n3252), .B(n3982), .Z(n3031) );
  HS65_LL_NOR2X6 U15499 ( .A(n3251), .B(n2917), .Z(n3636) );
  HS65_LL_NOR2X6 U15500 ( .A(n2883), .B(n2972), .Z(n3745) );
  HS65_LL_NOR2X6 U15501 ( .A(n2831), .B(n2997), .Z(n3860) );
  HS65_LL_NOR2X6 U15502 ( .A(n3095), .B(n2859), .Z(n3506) );
  HS65_LL_NOR2X6 U15503 ( .A(n3251), .B(n3047), .Z(n3552) );
  HS65_LL_NAND2X7 U15504 ( .A(n3197), .B(n2837), .Z(n3365) );
  HS65_LL_NAND2X7 U15505 ( .A(n2931), .B(n3116), .Z(n3080) );
  HS65_LL_NOR2X6 U15506 ( .A(n3252), .B(n3269), .Z(n3030) );
  HS65_LL_NOR2X6 U15507 ( .A(n8168), .B(n7724), .Z(n8821) );
  HS65_LL_NOR2X6 U15508 ( .A(n8145), .B(n7686), .Z(n8731) );
  HS65_LL_NOR2X6 U15509 ( .A(n3984), .B(n2917), .Z(n3283) );
  HS65_LL_NOR2X6 U15510 ( .A(n7660), .B(n7663), .Z(n8775) );
  HS65_LL_NOR2X6 U15511 ( .A(n7620), .B(n7623), .Z(n8685) );
  HS65_LL_NOR2X6 U15512 ( .A(n8057), .B(n8029), .Z(n8604) );
  HS65_LL_NOR2X6 U15513 ( .A(n2913), .B(n3034), .Z(n3027) );
  HS65_LL_NOR2X6 U15514 ( .A(n8168), .B(n8776), .Z(n7927) );
  HS65_LL_NOR2X6 U15515 ( .A(n8145), .B(n8686), .Z(n7829) );
  HS65_LL_NOR2X6 U15516 ( .A(n3928), .B(n2855), .Z(n3492) );
  HS65_LL_NOR2X6 U15517 ( .A(n3396), .B(n2846), .Z(n3181) );
  HS65_LL_NOR2X6 U15518 ( .A(n4747), .B(n4586), .Z(n5349) );
  HS65_LL_NOR2X6 U15519 ( .A(n4773), .B(n4603), .Z(n5464) );
  HS65_LL_NOR2X6 U15520 ( .A(n4627), .B(n4533), .Z(n5234) );
  HS65_LL_NOR2X6 U15521 ( .A(n6327), .B(n6179), .Z(n6941) );
  HS65_LL_NOR2X6 U15522 ( .A(n6366), .B(n6196), .Z(n7056) );
  HS65_LL_NOR2X6 U15523 ( .A(n6220), .B(n6126), .Z(n6826) );
  HS65_LL_NOR2X6 U15524 ( .A(n2995), .B(n3197), .Z(n3885) );
  HS65_LL_NOR2X6 U15525 ( .A(n2857), .B(n2931), .Z(n3531) );
  HS65_LL_NOR2X6 U15526 ( .A(n4566), .B(n4709), .Z(n5068) );
  HS65_LL_NOR2X6 U15527 ( .A(n6159), .B(n6302), .Z(n6661) );
  HS65_LL_NOR2X6 U15528 ( .A(n4734), .B(n4882), .Z(n5259) );
  HS65_LL_NOR2X6 U15529 ( .A(n4795), .B(n4994), .Z(n5374) );
  HS65_LL_NOR2X6 U15530 ( .A(n4649), .B(n4868), .Z(n5142) );
  HS65_LL_NOR2X6 U15531 ( .A(n6349), .B(n6475), .Z(n6851) );
  HS65_LL_NOR2X6 U15532 ( .A(n6388), .B(n6587), .Z(n6966) );
  HS65_LL_NOR2X6 U15533 ( .A(n6242), .B(n6461), .Z(n6734) );
  HS65_LL_NAND2X7 U15534 ( .A(n3034), .B(n3033), .Z(n3040) );
  HS65_LL_NOR2X6 U15535 ( .A(n4775), .B(n5554), .Z(n5413) );
  HS65_LL_NOR2X6 U15536 ( .A(n6368), .B(n7146), .Z(n7005) );
  HS65_LL_NOR2X6 U15537 ( .A(n4629), .B(n5579), .Z(n5182) );
  HS65_LL_NOR2X6 U15538 ( .A(n6222), .B(n7171), .Z(n6774) );
  HS65_LL_NOR2X6 U15539 ( .A(n6117), .B(n6402), .Z(n6435) );
  HS65_LL_NOR2X6 U15540 ( .A(n4524), .B(n4809), .Z(n4842) );
  HS65_LL_AOI212X4 U15541 ( .A(n646), .B(n3703), .C(n656), .D(n3704), .E(n3705), .Z(n3696) );
  HS65_LL_NAND2X7 U15542 ( .A(n2981), .B(n2882), .Z(n3704) );
  HS65_LL_NOR2X6 U15543 ( .A(n2913), .B(n3984), .Z(n3609) );
  HS65_LL_NAND2X7 U15544 ( .A(n6048), .B(n6515), .Z(n6346) );
  HS65_LL_NAND2X7 U15545 ( .A(n4494), .B(n4975), .Z(n4792) );
  HS65_LL_NAND2X7 U15546 ( .A(n4626), .B(n4847), .Z(n4646) );
  HS65_LL_NAND2X7 U15547 ( .A(n6219), .B(n6440), .Z(n6239) );
  HS65_LL_NAND2X7 U15548 ( .A(n4455), .B(n4922), .Z(n4730) );
  HS65_LL_NAND2X7 U15549 ( .A(n6087), .B(n6568), .Z(n6385) );
  HS65_LL_NOR2X6 U15550 ( .A(n7173), .B(n7170), .Z(n6743) );
  HS65_LL_NOR2X6 U15551 ( .A(n5581), .B(n5578), .Z(n5151) );
  HS65_LL_NOR2X6 U15552 ( .A(n5630), .B(n5629), .Z(n5383) );
  HS65_LL_NOR2X6 U15553 ( .A(n7222), .B(n7221), .Z(n6975) );
  HS65_LL_NOR2X6 U15554 ( .A(n4460), .B(n5532), .Z(n5283) );
  HS65_LL_NOR2X6 U15555 ( .A(n4499), .B(n5554), .Z(n5398) );
  HS65_LL_NOR2X6 U15556 ( .A(n4525), .B(n5579), .Z(n5166) );
  HS65_LL_NOR2X6 U15557 ( .A(n6053), .B(n7124), .Z(n6875) );
  HS65_LL_NOR2X6 U15558 ( .A(n6092), .B(n7146), .Z(n6990) );
  HS65_LL_NOR2X6 U15559 ( .A(n6118), .B(n7171), .Z(n6758) );
  HS65_LL_NOR2X6 U15560 ( .A(n2855), .B(n2933), .Z(n3093) );
  HS65_LL_NOR2X6 U15561 ( .A(n3114), .B(n3112), .Z(n2955) );
  HS65_LL_NOR2X6 U15562 ( .A(n7831), .B(n7620), .Z(n8412) );
  HS65_LL_NOR2X6 U15563 ( .A(n7870), .B(n7660), .Z(n8464) );
  HS65_LL_NOR4ABX2 U15564 ( .A(n3989), .B(n3990), .C(n3991), .D(n3992), .Z(
        n3908) );
  HS65_LL_OAI222X2 U15565 ( .A(n3984), .B(n3588), .C(n3982), .D(n2914), .E(
        n3035), .F(n3269), .Z(n3992) );
  HS65_LL_NOR3AX2 U15566 ( .A(n3243), .B(n3554), .C(n3031), .Z(n3989) );
  HS65_LL_OAI212X5 U15567 ( .A(n3575), .B(n3225), .C(n2915), .D(n3252), .E(
        n3993), .Z(n3991) );
  HS65_LL_NOR2X6 U15568 ( .A(n4710), .B(n4551), .Z(n5099) );
  HS65_LL_NOR2X6 U15569 ( .A(n6303), .B(n6144), .Z(n6692) );
  HS65_LL_NOR2X6 U15570 ( .A(n3047), .B(n3994), .Z(n3594) );
  HS65_LL_NOR2X6 U15571 ( .A(n5496), .B(n5572), .Z(n5213) );
  HS65_LL_NOR2X6 U15572 ( .A(n7088), .B(n7164), .Z(n6805) );
  HS65_LL_NOR2X6 U15573 ( .A(n7848), .B(n7960), .Z(n8100) );
  HS65_LL_NOR2X6 U15574 ( .A(n6127), .B(n7164), .Z(n6823) );
  HS65_LL_NOR2X6 U15575 ( .A(n4534), .B(n5572), .Z(n5231) );
  HS65_LL_NOR2X6 U15576 ( .A(n6305), .B(n6143), .Z(n6613) );
  HS65_LL_NOR2X6 U15577 ( .A(n4712), .B(n4550), .Z(n5020) );
  HS65_LL_NOR2X6 U15578 ( .A(n8178), .B(n7651), .Z(n8435) );
  HS65_LL_NOR2X6 U15579 ( .A(n8155), .B(n7631), .Z(n8383) );
  HS65_LL_NAND2X7 U15580 ( .A(n8169), .B(n8168), .Z(n7738) );
  HS65_LL_NAND2X7 U15581 ( .A(n8146), .B(n8145), .Z(n7700) );
  HS65_LL_NAND2X7 U15582 ( .A(n4550), .B(n4710), .Z(n4569) );
  HS65_LL_NAND2X7 U15583 ( .A(n6143), .B(n6303), .Z(n6162) );
  HS65_LL_NOR2X6 U15584 ( .A(n6160), .B(n7064), .Z(n6616) );
  HS65_LL_NOR2X6 U15585 ( .A(n4567), .B(n5472), .Z(n5023) );
  HS65_LL_NOR2X6 U15586 ( .A(n3588), .B(n3994), .Z(n3273) );
  HS65_LL_NAND2X7 U15587 ( .A(n2956), .B(n2856), .Z(n2929) );
  HS65_LL_NOR2X6 U15588 ( .A(n3380), .B(n3204), .Z(n3364) );
  HS65_LL_NOR2X6 U15589 ( .A(n7835), .B(n8145), .Z(n8695) );
  HS65_LL_NOR2X6 U15590 ( .A(n7874), .B(n8168), .Z(n8785) );
  HS65_LL_NOR2X6 U15591 ( .A(n8057), .B(n7942), .Z(n8056) );
  HS65_LL_NOR2X6 U15592 ( .A(n2992), .B(n3204), .Z(n3403) );
  HS65_LL_NOR2X6 U15593 ( .A(n3380), .B(n3193), .Z(n3795) );
  HS65_LL_NOR2X6 U15594 ( .A(n3096), .B(n2927), .Z(n3437) );
  HS65_LL_NOR2X6 U15595 ( .A(n7940), .B(n8540), .Z(n8570) );
  HS65_LL_NOR2X6 U15596 ( .A(n4566), .B(n5026), .Z(n5091) );
  HS65_LL_NOR2X6 U15597 ( .A(n6159), .B(n6619), .Z(n6684) );
  HS65_LL_NOR2X6 U15598 ( .A(n6241), .B(n6116), .Z(n6784) );
  HS65_LL_NOR2X6 U15599 ( .A(n4648), .B(n4523), .Z(n5192) );
  HS65_LL_NOR2X6 U15600 ( .A(n4478), .B(n4483), .Z(n4664) );
  HS65_LL_NOR2X6 U15601 ( .A(n6071), .B(n6076), .Z(n6257) );
  HS65_LL_NOR2X6 U15602 ( .A(n4747), .B(n4882), .Z(n5262) );
  HS65_LL_NOR2X6 U15603 ( .A(n4773), .B(n4994), .Z(n5377) );
  HS65_LL_NOR2X6 U15604 ( .A(n4627), .B(n4868), .Z(n5145) );
  HS65_LL_NOR2X6 U15605 ( .A(n6366), .B(n6587), .Z(n6969) );
  HS65_LL_NOR2X6 U15606 ( .A(n6220), .B(n6461), .Z(n6737) );
  HS65_LL_NOR2X6 U15607 ( .A(n6327), .B(n6475), .Z(n6854) );
  HS65_LL_NOR2X6 U15608 ( .A(n7094), .B(n7106), .Z(n6623) );
  HS65_LL_NOR2X6 U15609 ( .A(n5502), .B(n5514), .Z(n5030) );
  HS65_LL_NOR2X6 U15610 ( .A(n4670), .B(n5514), .Z(n5095) );
  HS65_LL_NOR2X6 U15611 ( .A(n6263), .B(n7106), .Z(n6688) );
  HS65_LL_NOR2X6 U15612 ( .A(n7163), .B(n6727), .Z(n6410) );
  HS65_LL_NOR2X6 U15613 ( .A(n5571), .B(n5135), .Z(n4817) );
  HS65_LL_NOR2X6 U15614 ( .A(n3252), .B(n3994), .Z(n3235) );
  HS65_LL_NOR2X6 U15615 ( .A(n3574), .B(n3042), .Z(n3249) );
  HS65_LL_NOR2X6 U15616 ( .A(n3326), .B(n3129), .Z(n3680) );
  HS65_LL_NOR2X6 U15617 ( .A(n2914), .B(n3994), .Z(n3650) );
  HS65_LL_NOR2X6 U15618 ( .A(n8173), .B(n7651), .Z(n8829) );
  HS65_LL_NOR2X6 U15619 ( .A(n8150), .B(n7631), .Z(n8739) );
  HS65_LL_CBI4I1X5 U15620 ( .A(n3061), .B(n2958), .C(n3475), .D(n3476), .Z(
        n3474) );
  HS65_LL_NOR2X6 U15621 ( .A(n7992), .B(n7961), .Z(n8219) );
  HS65_LL_NAND2X7 U15622 ( .A(n2884), .B(n2969), .Z(n3131) );
  HS65_LL_NOR2X6 U15623 ( .A(n7992), .B(n7860), .Z(n7988) );
  HS65_LL_NOR2X6 U15624 ( .A(n4566), .B(n4668), .Z(n4708) );
  HS65_LL_NOR2X6 U15625 ( .A(n6159), .B(n6261), .Z(n6301) );
  HS65_LL_CBI4I1X5 U15626 ( .A(n3032), .B(n2917), .C(n3280), .D(n3551), .Z(
        n4086) );
  HS65_LL_NOR2X6 U15627 ( .A(n3096), .B(n2939), .Z(n3079) );
  HS65_LL_NOR2X6 U15628 ( .A(n3464), .B(n2939), .Z(n3122) );
  HS65_LL_NOR2X6 U15629 ( .A(n3271), .B(n3574), .Z(n3570) );
  HS65_LL_NOR2X6 U15630 ( .A(n6088), .B(n7222), .Z(n6540) );
  HS65_LL_NOR2X6 U15631 ( .A(n6049), .B(n7180), .Z(n6487) );
  HS65_LL_NOR2X6 U15632 ( .A(n4456), .B(n5588), .Z(n4894) );
  HS65_LL_NOR2X6 U15633 ( .A(n4495), .B(n5630), .Z(n4947) );
  HS65_LL_NOR2X6 U15634 ( .A(n6441), .B(n7173), .Z(n6412) );
  HS65_LL_NOR2X6 U15635 ( .A(n4848), .B(n5581), .Z(n4819) );
  HS65_LL_CBI4I1X5 U15636 ( .A(n2884), .B(n2972), .C(n3293), .D(n3678), .Z(
        n4236) );
  HS65_LL_NOR2X6 U15637 ( .A(n5472), .B(n5508), .Z(n5107) );
  HS65_LL_NOR2X6 U15638 ( .A(n7874), .B(n7653), .Z(n8828) );
  HS65_LL_NOR2X6 U15639 ( .A(n7835), .B(n7633), .Z(n8738) );
  HS65_LL_NOR2X6 U15640 ( .A(n7064), .B(n7100), .Z(n6700) );
  HS65_LL_CBI4I1X5 U15641 ( .A(n7630), .B(n7686), .C(n7636), .D(n7687), .Z(
        n7685) );
  HS65_LL_CBI4I1X5 U15642 ( .A(n7650), .B(n7724), .C(n7657), .D(n7725), .Z(
        n7723) );
  HS65_LL_NOR2X6 U15643 ( .A(n7806), .B(n7633), .Z(n7793) );
  HS65_LL_NOR2X6 U15644 ( .A(n7869), .B(n7653), .Z(n7892) );
  HS65_LL_NOR2X6 U15645 ( .A(n2933), .B(n3475), .Z(n3508) );
  HS65_LL_NAND2X7 U15646 ( .A(n3032), .B(n2914), .Z(n3045) );
  HS65_LL_NOR2X6 U15647 ( .A(n7664), .B(n7656), .Z(n8800) );
  HS65_LL_NOR2X6 U15648 ( .A(n7624), .B(n7619), .Z(n8710) );
  HS65_LL_NAND2X7 U15649 ( .A(n4551), .B(n4549), .Z(n4561) );
  HS65_LL_NAND2X7 U15650 ( .A(n6144), .B(n6142), .Z(n6154) );
  HS65_LL_NOR2X6 U15651 ( .A(n7858), .B(n8238), .Z(n8269) );
  HS65_LL_NAND2X7 U15652 ( .A(n2146), .B(n1898), .Z(n1875) );
  HS65_LL_NOR2X6 U15653 ( .A(n3114), .B(n3095), .Z(n3119) );
  HS65_LL_NOR2X6 U15654 ( .A(n7751), .B(n8123), .Z(n8233) );
  HS65_LL_NOR2X6 U15655 ( .A(n7948), .B(n8049), .Z(n8609) );
  HS65_LL_NAND2X7 U15656 ( .A(n1770), .B(n1522), .Z(n1499) );
  HS65_LL_NAND2X7 U15657 ( .A(n2522), .B(n2274), .Z(n2251) );
  HS65_LL_NAND2X7 U15658 ( .A(n1394), .B(n1146), .Z(n1123) );
  HS65_LL_NOR2X6 U15659 ( .A(n2994), .B(n3185), .Z(n3791) );
  HS65_LL_NOR2X6 U15660 ( .A(n2856), .B(n2958), .Z(n3433) );
  HS65_LL_NOR2X6 U15661 ( .A(n3183), .B(n3412), .Z(n3842) );
  HS65_LL_NOR2X6 U15662 ( .A(n7980), .B(n8254), .Z(n8250) );
  HS65_LL_NAND4ABX3 U15663 ( .A(n5073), .B(n5074), .C(n5075), .D(n5076), .Z(
        n4543) );
  HS65_LL_AOI212X4 U15664 ( .A(n45), .B(n5077), .C(n34), .D(n5078), .E(n5079), 
        .Z(n5076) );
  HS65_LL_AOI222X2 U15665 ( .A(n39), .B(n14), .C(n18), .D(n31), .E(n15), .F(
        n40), .Z(n5075) );
  HS65_LL_MX41X7 U15666 ( .D0(n24), .S0(n47), .D1(n20), .S1(n30), .D2(n37), 
        .S2(n4481), .D3(n42), .S3(n22), .Z(n5073) );
  HS65_LL_NAND4ABX3 U15667 ( .A(n6666), .B(n6667), .C(n6668), .D(n6669), .Z(
        n6136) );
  HS65_LL_AOI212X4 U15668 ( .A(n567), .B(n6670), .C(n556), .D(n6671), .E(n6672), .Z(n6669) );
  HS65_LL_AOI222X2 U15669 ( .A(n561), .B(n536), .C(n540), .D(n553), .E(n537), 
        .F(n562), .Z(n6668) );
  HS65_LL_MX41X7 U15670 ( .D0(n546), .S0(n569), .D1(n542), .S1(n552), .D2(n559), .S2(n6074), .D3(n564), .S3(n544), .Z(n6666) );
  HS65_LL_NAND4ABX3 U15671 ( .A(n5311), .B(n5312), .C(n5313), .D(n5314), .Z(
        n4741) );
  HS65_LL_AOI212X4 U15672 ( .A(n253), .B(n5315), .C(n263), .D(n5316), .E(n5317), .Z(n5314) );
  HS65_LL_NAND4ABX3 U15673 ( .A(n5318), .B(n5319), .C(n5320), .D(n5321), .Z(
        n5312) );
  HS65_LL_MX41X7 U15674 ( .D0(n234), .S0(n252), .D1(n238), .S1(n259), .D2(n261), .S2(n4589), .D3(n264), .S3(n232), .Z(n5311) );
  HS65_LL_NAND4ABX3 U15675 ( .A(n5426), .B(n5427), .C(n5428), .D(n5429), .Z(
        n4767) );
  HS65_LL_AOI212X4 U15676 ( .A(n470), .B(n5430), .C(n480), .D(n5431), .E(n5432), .Z(n5429) );
  HS65_LL_NAND4ABX3 U15677 ( .A(n5433), .B(n5434), .C(n5435), .D(n5436), .Z(
        n5427) );
  HS65_LL_MX41X7 U15678 ( .D0(n451), .S0(n469), .D1(n455), .S1(n476), .D2(n478), .S2(n4606), .D3(n481), .S3(n449), .Z(n5426) );
  HS65_LL_NAND4ABX3 U15679 ( .A(n6903), .B(n6904), .C(n6905), .D(n6906), .Z(
        n6321) );
  HS65_LL_AOI212X4 U15680 ( .A(n88), .B(n6907), .C(n86), .D(n6908), .E(n6909), 
        .Z(n6906) );
  HS65_LL_NAND4ABX3 U15681 ( .A(n6910), .B(n6911), .C(n6912), .D(n6913), .Z(
        n6904) );
  HS65_LL_MX41X7 U15682 ( .D0(n63), .S0(n89), .D1(n60), .S1(n77), .D2(n85), 
        .S2(n6182), .D3(n78), .S3(n65), .Z(n6903) );
  HS65_LL_NAND4ABX3 U15683 ( .A(n5195), .B(n5196), .C(n5197), .D(n5198), .Z(
        n4620) );
  HS65_LL_AOI212X4 U15684 ( .A(n700), .B(n5199), .C(n689), .D(n5200), .E(n5201), .Z(n5198) );
  HS65_LL_NAND4ABX3 U15685 ( .A(n5202), .B(n5203), .C(n5204), .D(n5205), .Z(
        n5196) );
  HS65_LL_MX41X7 U15686 ( .D0(n679), .S0(n702), .D1(n675), .S1(n685), .D2(n692), .S2(n4521), .D3(n697), .S3(n677), .Z(n5195) );
  HS65_LL_NAND4ABX3 U15687 ( .A(n7018), .B(n7019), .C(n7020), .D(n7021), .Z(
        n6360) );
  HS65_LL_AOI212X4 U15688 ( .A(n295), .B(n7022), .C(n305), .D(n7023), .E(n7024), .Z(n7021) );
  HS65_LL_NAND4ABX3 U15689 ( .A(n7025), .B(n7026), .C(n7027), .D(n7028), .Z(
        n7019) );
  HS65_LL_MX41X7 U15690 ( .D0(n276), .S0(n294), .D1(n280), .S1(n301), .D2(n303), .S2(n6199), .D3(n306), .S3(n274), .Z(n7018) );
  HS65_LL_NAND4ABX3 U15691 ( .A(n6787), .B(n6788), .C(n6789), .D(n6790), .Z(
        n6213) );
  HS65_LL_AOI212X4 U15692 ( .A(n524), .B(n6791), .C(n513), .D(n6792), .E(n6793), .Z(n6790) );
  HS65_LL_NAND4ABX3 U15693 ( .A(n6794), .B(n6795), .C(n6796), .D(n6797), .Z(
        n6788) );
  HS65_LL_MX41X7 U15694 ( .D0(n503), .S0(n526), .D1(n499), .S1(n509), .D2(n516), .S2(n6114), .D3(n521), .S3(n501), .Z(n6787) );
  HS65_LL_NOR2X6 U15695 ( .A(n3286), .B(n3280), .Z(n3567) );
  HS65_LL_NOR2X6 U15696 ( .A(n2969), .B(n3158), .Z(n3676) );
  HS65_LL_NOR2X6 U15697 ( .A(n7099), .B(n6606), .Z(n6272) );
  HS65_LL_NOR2X6 U15698 ( .A(n5507), .B(n5013), .Z(n4679) );
  HS65_LL_NOR2X6 U15699 ( .A(n7806), .B(n7623), .Z(n8154) );
  HS65_LL_NOR2X6 U15700 ( .A(n7869), .B(n7663), .Z(n8177) );
  HS65_LL_NOR2X6 U15701 ( .A(n1609), .B(n1545), .Z(n1593) );
  HS65_LL_NOR2X6 U15702 ( .A(n5265), .B(n4923), .Z(n4750) );
  HS65_LL_NOR2X6 U15703 ( .A(n5380), .B(n4976), .Z(n4777) );
  HS65_LL_NOR2X6 U15704 ( .A(n5148), .B(n4849), .Z(n4631) );
  HS65_LL_NOR2X6 U15705 ( .A(n6857), .B(n6516), .Z(n6331) );
  HS65_LL_NOR2X6 U15706 ( .A(n6972), .B(n6569), .Z(n6370) );
  HS65_LL_NOR2X6 U15707 ( .A(n6740), .B(n6442), .Z(n6224) );
  HS65_LL_NOR2X6 U15708 ( .A(n6302), .B(n7094), .Z(n6273) );
  HS65_LL_NOR2X6 U15709 ( .A(n4709), .B(n5502), .Z(n4680) );
  HS65_LL_NOR2X6 U15710 ( .A(n3286), .B(n3224), .Z(n3651) );
  HS65_LL_NOR2X6 U15711 ( .A(n8048), .B(n8556), .Z(n8553) );
  HS65_LL_NOR2X6 U15712 ( .A(n3286), .B(n3043), .Z(n3635) );
  HS65_LL_NOR2X6 U15713 ( .A(n4485), .B(n4572), .Z(n5050) );
  HS65_LL_NOR2X6 U15714 ( .A(n6078), .B(n6165), .Z(n6643) );
  HS65_LL_AOI12X2 U15715 ( .A(n6076), .B(n6077), .C(n6078), .Z(n6075) );
  HS65_LL_AOI12X2 U15716 ( .A(n4483), .B(n4484), .C(n4485), .Z(n4482) );
  HS65_LL_NOR2X6 U15717 ( .A(n3252), .B(n3043), .Z(n3554) );
  HS65_LL_NOR2X6 U15718 ( .A(n2914), .B(n3054), .Z(n3557) );
  HS65_LL_NOR2X6 U15719 ( .A(n8313), .B(n7952), .Z(n8366) );
  HS65_LL_NOR2X6 U15720 ( .A(n3033), .B(n3271), .Z(n3637) );
  HS65_LL_NOR2X6 U15721 ( .A(n8155), .B(n7619), .Z(n8153) );
  HS65_LL_NOR2X6 U15722 ( .A(n8178), .B(n7656), .Z(n8176) );
  HS65_LL_NAND2X7 U15723 ( .A(n4484), .B(n4668), .Z(n5478) );
  HS65_LL_NAND2X7 U15724 ( .A(n6077), .B(n6261), .Z(n7070) );
  HS65_LL_NOR2X6 U15725 ( .A(n2918), .B(n3574), .Z(n3561) );
  HS65_LL_NOR4ABX2 U15726 ( .A(n8141), .B(n8142), .C(n8143), .D(n8144), .Z(
        n8000) );
  HS65_LL_NOR3X4 U15727 ( .A(n7673), .B(n8153), .C(n8154), .Z(n8141) );
  HS65_LL_OAI212X5 U15728 ( .A(n7630), .B(n8145), .C(n8146), .D(n7624), .E(
        n8147), .Z(n8144) );
  HS65_LL_NAND3AX6 U15729 ( .A(n7812), .B(n8148), .C(n8149), .Z(n8143) );
  HS65_LL_NOR4ABX2 U15730 ( .A(n8164), .B(n8165), .C(n8166), .D(n8167), .Z(
        n8013) );
  HS65_LL_NOR3X4 U15731 ( .A(n7711), .B(n8176), .C(n8177), .Z(n8164) );
  HS65_LL_OAI212X5 U15732 ( .A(n7650), .B(n8168), .C(n8169), .D(n7664), .E(
        n8170), .Z(n8167) );
  HS65_LL_NAND3AX6 U15733 ( .A(n7910), .B(n8171), .C(n8172), .Z(n8166) );
  HS65_LL_NOR2X6 U15734 ( .A(n4975), .B(n4774), .Z(n5465) );
  HS65_LL_NOR2X6 U15735 ( .A(n4922), .B(n4748), .Z(n5350) );
  HS65_LL_NOR2X6 U15736 ( .A(n6568), .B(n6367), .Z(n7057) );
  HS65_LL_NOR2X6 U15737 ( .A(n4847), .B(n4628), .Z(n5235) );
  HS65_LL_NOR2X6 U15738 ( .A(n6440), .B(n6221), .Z(n6827) );
  HS65_LL_NOR2X6 U15739 ( .A(n6515), .B(n6328), .Z(n6942) );
  HS65_LL_NOR2X6 U15740 ( .A(n4868), .B(n4523), .Z(n5186) );
  HS65_LL_NOR2X6 U15741 ( .A(n6461), .B(n6116), .Z(n6778) );
  HS65_LL_NOR2X6 U15742 ( .A(n8057), .B(n8039), .Z(n8323) );
  HS65_LL_NOR2X6 U15743 ( .A(n5554), .B(n4976), .Z(n4783) );
  HS65_LL_NOR2X6 U15744 ( .A(n5579), .B(n4849), .Z(n4637) );
  HS65_LL_NOR2X6 U15745 ( .A(n7171), .B(n6442), .Z(n6230) );
  HS65_LL_NOR2X6 U15746 ( .A(n7146), .B(n6569), .Z(n6376) );
  HS65_LL_NOR2X6 U15747 ( .A(n5532), .B(n4923), .Z(n4756) );
  HS65_LL_NOR2X6 U15748 ( .A(n7124), .B(n6516), .Z(n6337) );
  HS65_LL_NOR2X6 U15749 ( .A(n8155), .B(n7822), .Z(n7673) );
  HS65_LL_NOR2X6 U15750 ( .A(n8178), .B(n7920), .Z(n7711) );
  HS65_LL_NOR4ABX2 U15751 ( .A(n6138), .B(n6139), .C(n6140), .D(n6141), .Z(
        n6067) );
  HS65_LL_NAND4ABX3 U15752 ( .A(n6147), .B(n6148), .C(n6149), .D(n6150), .Z(
        n6140) );
  HS65_LL_NOR3AX2 U15753 ( .A(n6155), .B(n6156), .C(n6157), .Z(n6138) );
  HS65_LL_OAI212X5 U15754 ( .A(n6142), .B(n6143), .C(n6144), .D(n6145), .E(
        n6146), .Z(n6141) );
  HS65_LL_NOR4ABX2 U15755 ( .A(n4545), .B(n4546), .C(n4547), .D(n4548), .Z(
        n4474) );
  HS65_LL_NAND4ABX3 U15756 ( .A(n4554), .B(n4555), .C(n4556), .D(n4557), .Z(
        n4547) );
  HS65_LL_NOR3AX2 U15757 ( .A(n4562), .B(n4563), .C(n4564), .Z(n4545) );
  HS65_LL_OAI212X5 U15758 ( .A(n4549), .B(n4550), .C(n4551), .D(n4552), .E(
        n4553), .Z(n4548) );
  HS65_LL_NAND2X7 U15759 ( .A(n3972), .B(n2995), .Z(n2843) );
  HS65_LL_NOR2X6 U15760 ( .A(n3588), .B(n3224), .Z(n3632) );
  HS65_LL_NOR2X6 U15761 ( .A(n4789), .B(n4995), .Z(n4974) );
  HS65_LL_NOR2X6 U15762 ( .A(n4727), .B(n4883), .Z(n4921) );
  HS65_LL_NOR2X6 U15763 ( .A(n6382), .B(n6588), .Z(n6567) );
  HS65_LL_NOR2X6 U15764 ( .A(n6343), .B(n6476), .Z(n6514) );
  HS65_LL_NOR2X6 U15765 ( .A(n6236), .B(n6462), .Z(n6439) );
  HS65_LL_NOR2X6 U15766 ( .A(n4643), .B(n4869), .Z(n4846) );
  HS65_LL_NOR2X6 U15767 ( .A(n3097), .B(n3067), .Z(n3470) );
  HS65_LL_NOR2X6 U15768 ( .A(n5267), .B(n5591), .Z(n5317) );
  HS65_LL_NOR2X6 U15769 ( .A(n5382), .B(n5616), .Z(n5432) );
  HS65_LL_NOR2X6 U15770 ( .A(n6859), .B(n7183), .Z(n6909) );
  HS65_LL_NOR2X6 U15771 ( .A(n5150), .B(n5572), .Z(n5201) );
  HS65_LL_NOR2X6 U15772 ( .A(n6974), .B(n7208), .Z(n7024) );
  HS65_LL_NOR2X6 U15773 ( .A(n6742), .B(n7164), .Z(n6793) );
  HS65_LL_NOR2X6 U15774 ( .A(n2956), .B(n3097), .Z(n3486) );
  HS65_LL_NOR2X6 U15775 ( .A(n2832), .B(n2829), .Z(n3841) );
  HS65_LL_NAND4ABX3 U15776 ( .A(n3681), .B(n3682), .C(n3683), .D(n3684), .Z(
        n3302) );
  HS65_LL_AOI222X2 U15777 ( .A(n658), .B(n638), .C(n650), .D(n3131), .E(n640), 
        .F(n651), .Z(n3683) );
  HS65_LL_OAI212X5 U15778 ( .A(n3691), .B(n3692), .C(n3693), .D(n3342), .E(
        n3694), .Z(n3681) );
  HS65_LL_NAND4ABX3 U15779 ( .A(n3688), .B(n2892), .C(n3689), .D(n3690), .Z(
        n3682) );
  HS65_LL_NOR4ABX2 U15780 ( .A(n4743), .B(n4744), .C(n4745), .D(n4746), .Z(
        n4583) );
  HS65_LL_NOR3X4 U15781 ( .A(n4758), .B(n4759), .C(n4760), .Z(n4743) );
  HS65_LL_OAI212X5 U15782 ( .A(n4455), .B(n4747), .C(n4748), .D(n4733), .E(
        n4749), .Z(n4746) );
  HS65_LL_NAND4ABX3 U15783 ( .A(n4750), .B(n4751), .C(n4752), .D(n4753), .Z(
        n4745) );
  HS65_LL_NOR4ABX2 U15784 ( .A(n6215), .B(n6216), .C(n6217), .D(n6218), .Z(
        n6123) );
  HS65_LL_NOR3X4 U15785 ( .A(n6232), .B(n6233), .C(n6234), .Z(n6215) );
  HS65_LL_OAI212X5 U15786 ( .A(n6219), .B(n6220), .C(n6221), .D(n6222), .E(
        n6223), .Z(n6218) );
  HS65_LL_NAND4ABX3 U15787 ( .A(n6224), .B(n6225), .C(n6226), .D(n6227), .Z(
        n6217) );
  HS65_LL_NOR4ABX2 U15788 ( .A(n4769), .B(n4770), .C(n4771), .D(n4772), .Z(
        n4600) );
  HS65_LL_NOR3X4 U15789 ( .A(n4785), .B(n4786), .C(n4787), .Z(n4769) );
  HS65_LL_OAI212X5 U15790 ( .A(n4494), .B(n4773), .C(n4774), .D(n4775), .E(
        n4776), .Z(n4772) );
  HS65_LL_NAND4ABX3 U15791 ( .A(n4777), .B(n4778), .C(n4779), .D(n4780), .Z(
        n4771) );
  HS65_LL_NOR4ABX2 U15792 ( .A(n6362), .B(n6363), .C(n6364), .D(n6365), .Z(
        n6193) );
  HS65_LL_NOR3X4 U15793 ( .A(n6378), .B(n6379), .C(n6380), .Z(n6362) );
  HS65_LL_OAI212X5 U15794 ( .A(n6087), .B(n6366), .C(n6367), .D(n6368), .E(
        n6369), .Z(n6365) );
  HS65_LL_NAND4ABX3 U15795 ( .A(n6370), .B(n6371), .C(n6372), .D(n6373), .Z(
        n6364) );
  HS65_LL_NOR4ABX2 U15796 ( .A(n6323), .B(n6324), .C(n6325), .D(n6326), .Z(
        n6176) );
  HS65_LL_NOR3X4 U15797 ( .A(n6339), .B(n6340), .C(n6341), .Z(n6323) );
  HS65_LL_OAI212X5 U15798 ( .A(n6048), .B(n6327), .C(n6328), .D(n6329), .E(
        n6330), .Z(n6326) );
  HS65_LL_NAND4ABX3 U15799 ( .A(n6331), .B(n6332), .C(n6333), .D(n6334), .Z(
        n6325) );
  HS65_LL_NOR4ABX2 U15800 ( .A(n4622), .B(n4623), .C(n4624), .D(n4625), .Z(
        n4530) );
  HS65_LL_NOR3X4 U15801 ( .A(n4639), .B(n4640), .C(n4641), .Z(n4622) );
  HS65_LL_OAI212X5 U15802 ( .A(n4626), .B(n4627), .C(n4628), .D(n4629), .E(
        n4630), .Z(n4625) );
  HS65_LL_NAND4ABX3 U15803 ( .A(n4631), .B(n4632), .C(n4633), .D(n4634), .Z(
        n4624) );
  HS65_LL_NOR2X6 U15804 ( .A(n7851), .B(n8649), .Z(n7984) );
  HS65_LL_NOR2AX3 U15805 ( .A(n4521), .B(n4524), .Z(n5143) );
  HS65_LL_NOR2AX3 U15806 ( .A(n6114), .B(n6117), .Z(n6735) );
  HS65_LL_NAND2X7 U15807 ( .A(n3807), .B(n2995), .Z(n3384) );
  HS65_LL_NOR2X6 U15808 ( .A(n4549), .B(n4670), .Z(n4707) );
  HS65_LL_NOR2X6 U15809 ( .A(n6142), .B(n6263), .Z(n6300) );
  HS65_LL_NOR2X6 U15810 ( .A(n3491), .B(n2938), .Z(n3493) );
  HS65_LL_NOR2X6 U15811 ( .A(n3116), .B(n2938), .Z(n3509) );
  HS65_LL_NOR2X6 U15812 ( .A(n4567), .B(n4670), .Z(n5044) );
  HS65_LL_NOR2X6 U15813 ( .A(n6160), .B(n6263), .Z(n6637) );
  HS65_LL_NAND2X7 U15814 ( .A(n3952), .B(n2970), .Z(n2895) );
  HS65_LL_NOR2X6 U15815 ( .A(n7662), .B(n8173), .Z(n7710) );
  HS65_LL_NOR2X6 U15816 ( .A(n7633), .B(n7620), .Z(n8750) );
  HS65_LL_NOR2X6 U15817 ( .A(n7653), .B(n7660), .Z(n8840) );
  HS65_LL_NAND2X7 U15818 ( .A(n4093), .B(n2915), .Z(n3912) );
  HS65_LL_NAND2X7 U15819 ( .A(n3928), .B(n2857), .Z(n3897) );
  HS65_LL_NOR2X6 U15820 ( .A(n5501), .B(n4711), .Z(n4560) );
  HS65_LL_NOR2X6 U15821 ( .A(n7093), .B(n6304), .Z(n6153) );
  HS65_LL_NOR2X6 U15822 ( .A(n7650), .B(n7714), .Z(n7888) );
  HS65_LL_NOR2X6 U15823 ( .A(n3252), .B(n4093), .Z(n3258) );
  HS65_LL_NOR2X6 U15824 ( .A(n8049), .B(n7767), .Z(n8345) );
  HS65_LL_NOR2X6 U15825 ( .A(n3183), .B(n2994), .Z(n3801) );
  HS65_LL_NAND2X7 U15826 ( .A(n3047), .B(n3271), .Z(n3236) );
  HS65_LL_NOR2X6 U15827 ( .A(n3157), .B(n3731), .Z(n3728) );
  HS65_LL_NOR2X6 U15828 ( .A(n6085), .B(n6587), .Z(n6958) );
  HS65_LL_NOR2X6 U15829 ( .A(n4850), .B(n4868), .Z(n5133) );
  HS65_LL_NOR2X6 U15830 ( .A(n6443), .B(n6461), .Z(n6725) );
  HS65_LL_NOR2X6 U15831 ( .A(n6046), .B(n6475), .Z(n6843) );
  HS65_LL_NOR2X6 U15832 ( .A(n4453), .B(n4882), .Z(n5251) );
  HS65_LL_NOR2X6 U15833 ( .A(n4492), .B(n4994), .Z(n5366) );
  HS65_LL_IVX9 U15834 ( .A(n8686), .Z(n593) );
  HS65_LL_CBI4I1X5 U15835 ( .A(n3280), .B(n3034), .C(n3053), .D(n3600), .Z(
        n3599) );
  HS65_LL_NOR2X6 U15836 ( .A(n7981), .B(n7749), .Z(n8112) );
  HS65_LL_NOR2X6 U15837 ( .A(n8527), .B(n7941), .Z(n8522) );
  HS65_LL_NAND2X7 U15838 ( .A(n8005), .B(n8421), .Z(n7841) );
  HS65_LL_NAND2X7 U15839 ( .A(n8018), .B(n8473), .Z(n7880) );
  HS65_LL_NOR2X6 U15840 ( .A(n3157), .B(n2969), .Z(n3686) );
  HS65_LL_NOR2X6 U15841 ( .A(n3042), .B(n2915), .Z(n3250) );
  HS65_LL_NOR2X6 U15842 ( .A(n3183), .B(n2845), .Z(n3379) );
  HS65_LL_NOR2X6 U15843 ( .A(n3157), .B(n2875), .Z(n3325) );
  HS65_LL_NOR2X6 U15844 ( .A(n8048), .B(n7767), .Z(n8338) );
  HS65_LL_NAND2X7 U15845 ( .A(n3270), .B(n3271), .Z(n3585) );
  HS65_LL_NOR4ABX2 U15846 ( .A(n5631), .B(n5632), .C(n5633), .D(n5634), .Z(
        n5543) );
  HS65_LL_OAI222X2 U15847 ( .A(n4610), .B(n5629), .C(n5554), .D(n4975), .E(
        n5380), .F(n4775), .Z(n5634) );
  HS65_LL_NOR3X4 U15848 ( .A(n4783), .B(n5410), .C(n5454), .Z(n5631) );
  HS65_LL_OAI212X5 U15849 ( .A(n5449), .B(n4509), .C(n4976), .D(n4995), .E(
        n5635), .Z(n5633) );
  HS65_LL_NOR4ABX2 U15850 ( .A(n5574), .B(n5575), .C(n5576), .D(n5577), .Z(
        n5487) );
  HS65_LL_OAI222X2 U15851 ( .A(n5135), .B(n5578), .C(n5579), .D(n4847), .E(
        n5148), .F(n4629), .Z(n5577) );
  HS65_LL_NOR3X4 U15852 ( .A(n4637), .B(n5179), .C(n5224), .Z(n5574) );
  HS65_LL_OAI212X5 U15853 ( .A(n5219), .B(n4809), .C(n4849), .D(n4869), .E(
        n5580), .Z(n5576) );
  HS65_LL_NOR4ABX2 U15854 ( .A(n7166), .B(n7167), .C(n7168), .D(n7169), .Z(
        n7079) );
  HS65_LL_OAI222X2 U15855 ( .A(n6727), .B(n7170), .C(n7171), .D(n6440), .E(
        n6740), .F(n6222), .Z(n7169) );
  HS65_LL_NOR3X4 U15856 ( .A(n6230), .B(n6771), .C(n6816), .Z(n7166) );
  HS65_LL_OAI212X5 U15857 ( .A(n6811), .B(n6402), .C(n6442), .D(n6462), .E(
        n7172), .Z(n7168) );
  HS65_LL_NOR4ABX2 U15858 ( .A(n7223), .B(n7224), .C(n7225), .D(n7226), .Z(
        n7135) );
  HS65_LL_OAI222X2 U15859 ( .A(n6203), .B(n7221), .C(n7146), .D(n6568), .E(
        n6972), .F(n6368), .Z(n7226) );
  HS65_LL_NOR3X4 U15860 ( .A(n6376), .B(n7002), .C(n7046), .Z(n7223) );
  HS65_LL_OAI212X5 U15861 ( .A(n7041), .B(n6102), .C(n6569), .D(n6588), .E(
        n7227), .Z(n7225) );
  HS65_LL_NOR4ABX2 U15862 ( .A(n5605), .B(n5606), .C(n5607), .D(n5608), .Z(
        n5521) );
  HS65_LL_OAI222X2 U15863 ( .A(n4593), .B(n5604), .C(n5532), .D(n4922), .E(
        n5265), .F(n4733), .Z(n5608) );
  HS65_LL_NOR3X4 U15864 ( .A(n4756), .B(n5295), .C(n5339), .Z(n5605) );
  HS65_LL_OAI212X5 U15865 ( .A(n5334), .B(n4448), .C(n4923), .D(n4883), .E(
        n5609), .Z(n5607) );
  HS65_LL_CBI4I1X5 U15866 ( .A(n7636), .B(n8146), .C(n7632), .D(n8676), .Z(
        n8675) );
  HS65_LL_CBI4I1X5 U15867 ( .A(n7657), .B(n8169), .C(n7652), .D(n8766), .Z(
        n8765) );
  HS65_LL_NAND2X7 U15868 ( .A(n3692), .B(n2970), .Z(n3330) );
  HS65_LL_NOR2X6 U15869 ( .A(n3615), .B(n3982), .Z(n3617) );
  HS65_LL_NOR2X6 U15870 ( .A(n3380), .B(n2831), .Z(n3402) );
  HS65_LL_NOR2X6 U15871 ( .A(n2958), .B(n3067), .Z(n2954) );
  HS65_LL_NOR2X6 U15872 ( .A(n2957), .B(n3096), .Z(n3432) );
  HS65_LL_NAND2X7 U15873 ( .A(n5630), .B(n4500), .Z(n5430) );
  HS65_LL_NAND2X7 U15874 ( .A(n7222), .B(n6093), .Z(n7022) );
  HS65_LL_NAND2X7 U15875 ( .A(n5581), .B(n5496), .Z(n5199) );
  HS65_LL_NAND2X7 U15876 ( .A(n7173), .B(n7088), .Z(n6791) );
  HS65_LL_NOR2X6 U15877 ( .A(n5028), .B(n5508), .Z(n5079) );
  HS65_LL_NOR2X6 U15878 ( .A(n6621), .B(n7100), .Z(n6672) );
  HS65_LL_NOR2X6 U15879 ( .A(n3846), .B(n3406), .Z(n3363) );
  HS65_LL_NOR2X6 U15880 ( .A(n3193), .B(n3412), .Z(n2839) );
  HS65_LL_NOR2X6 U15881 ( .A(n2927), .B(n3067), .Z(n3503) );
  HS65_LL_NOR4ABX2 U15882 ( .A(n8972), .B(n8973), .C(n8974), .D(n8975), .Z(
        n8483) );
  HS65_LL_OAI222X2 U15883 ( .A(n8649), .B(n8207), .C(n7860), .D(n7847), .E(
        n7993), .F(n7966), .Z(n8975) );
  HS65_LL_NOR3X4 U15884 ( .A(n7988), .B(n8284), .C(n8219), .Z(n8972) );
  HS65_LL_OAI212X5 U15885 ( .A(n8303), .B(n7749), .C(n7848), .D(n7992), .E(
        n8976), .Z(n8974) );
  HS65_LL_NOR4ABX2 U15886 ( .A(n4037), .B(n4038), .C(n4039), .D(n4040), .Z(
        n3957) );
  HS65_LL_OAI222X2 U15887 ( .A(n3970), .B(n2992), .C(n3203), .D(n2994), .E(
        n3397), .F(n3184), .Z(n4040) );
  HS65_LL_NOR3X4 U15888 ( .A(n3795), .B(n3187), .C(n3381), .Z(n4037) );
  HS65_LL_NOR4ABX2 U15889 ( .A(n3849), .B(n3411), .C(n3877), .D(n3860), .Z(
        n4038) );
  HS65_LL_NOR2X6 U15890 ( .A(n3326), .B(n2883), .Z(n3348) );
  HS65_LL_NOR2X6 U15891 ( .A(n3069), .B(n2855), .Z(n3098) );
  HS65_LL_NOR2X6 U15892 ( .A(n8313), .B(n8510), .Z(n7764) );
  HS65_LL_NOR2X6 U15893 ( .A(n3096), .B(n3095), .Z(n3121) );
  HS65_LL_NOR2X6 U15894 ( .A(n3129), .B(n3299), .Z(n2891) );
  HS65_LL_NOR4ABX2 U15895 ( .A(n3922), .B(n3923), .C(n3924), .D(n3925), .Z(
        n3893) );
  HS65_LL_OAI222X2 U15896 ( .A(n3926), .B(n3464), .C(n2938), .D(n2856), .E(
        n3115), .F(n2932), .Z(n3925) );
  HS65_LL_NOR3X4 U15897 ( .A(n3437), .B(n2960), .C(n3098), .Z(n3922) );
  HS65_LL_NOR4ABX2 U15898 ( .A(n3494), .B(n3066), .C(n3523), .D(n3506), .Z(
        n3923) );
  HS65_LL_NOR4ABX2 U15899 ( .A(n5510), .B(n5511), .C(n5512), .D(n5513), .Z(
        n5473) );
  HS65_LL_OAI222X2 U15900 ( .A(n5013), .B(n5514), .C(n5501), .D(n4710), .E(
        n5026), .F(n4552), .Z(n5513) );
  HS65_LL_NOR3X4 U15901 ( .A(n4560), .B(n5057), .C(n5088), .Z(n5510) );
  HS65_LL_OAI212X5 U15902 ( .A(n5113), .B(n4670), .C(n4711), .D(n4668), .E(
        n5515), .Z(n5512) );
  HS65_LL_NOR4ABX2 U15903 ( .A(n7102), .B(n7103), .C(n7104), .D(n7105), .Z(
        n7065) );
  HS65_LL_OAI222X2 U15904 ( .A(n6606), .B(n7106), .C(n7093), .D(n6303), .E(
        n6619), .F(n6145), .Z(n7105) );
  HS65_LL_NOR3X4 U15905 ( .A(n6153), .B(n6650), .C(n6681), .Z(n7102) );
  HS65_LL_OAI212X5 U15906 ( .A(n6706), .B(n6263), .C(n6304), .D(n6261), .E(
        n7107), .Z(n7104) );
  HS65_LL_NOR2X6 U15907 ( .A(n4567), .B(n4667), .Z(n5048) );
  HS65_LL_NOR2X6 U15908 ( .A(n6160), .B(n6260), .Z(n6641) );
  HS65_LL_NOR2X6 U15909 ( .A(n2830), .B(n3807), .Z(n3790) );
  HS65_LL_NOR2X6 U15910 ( .A(n3185), .B(n3412), .Z(n3182) );
  HS65_LL_NOR2X6 U15911 ( .A(n4712), .B(n4667), .Z(n5011) );
  HS65_LL_NOR2X6 U15912 ( .A(n6305), .B(n6260), .Z(n6604) );
  HS65_LL_NOR4ABX2 U15913 ( .A(n8920), .B(n8921), .C(n8922), .D(n8923), .Z(
        n8849) );
  HS65_LL_OAI222X2 U15914 ( .A(n8630), .B(n8510), .C(n7942), .D(n7948), .E(
        n8058), .F(n8034), .Z(n8923) );
  HS65_LL_NOR3X4 U15915 ( .A(n8056), .B(n8583), .C(n8604), .Z(n8920) );
  HS65_LL_OAI212X5 U15916 ( .A(n8528), .B(n7767), .C(n7949), .D(n8057), .E(
        n8927), .Z(n8922) );
  HS65_LL_NOR2X6 U15917 ( .A(n3984), .B(n3286), .Z(n3649) );
  HS65_LL_NAND2X7 U15918 ( .A(n4608), .B(n4995), .Z(n4506) );
  HS65_LL_NAND2X7 U15919 ( .A(n4591), .B(n4883), .Z(n4467) );
  HS65_LL_NAND2X7 U15920 ( .A(n4524), .B(n4869), .Z(n5492) );
  HS65_LL_NAND2X7 U15921 ( .A(n6201), .B(n6588), .Z(n6099) );
  HS65_LL_NAND2X7 U15922 ( .A(n6117), .B(n6462), .Z(n7084) );
  HS65_LL_NAND2X7 U15923 ( .A(n6184), .B(n6476), .Z(n6060) );
  HS65_LL_NOR2X6 U15924 ( .A(n3269), .B(n3053), .Z(n3582) );
  HS65_LL_NAND2X7 U15925 ( .A(n2832), .B(n2994), .Z(n3195) );
  HS65_LL_NOR2X6 U15926 ( .A(n7768), .B(n8630), .Z(n8557) );
  HS65_LL_NOR2X6 U15927 ( .A(n7952), .B(n8630), .Z(n8052) );
  HS65_LL_NOR2X6 U15928 ( .A(n3491), .B(n3061), .Z(n3078) );
  HS65_LL_NOR4ABX2 U15929 ( .A(n9087), .B(n9088), .C(n9089), .D(n9090), .Z(
        n7646) );
  HS65_LL_OAI222X2 U15930 ( .A(n7663), .B(n7919), .C(n7656), .D(n8449), .E(
        n7664), .F(n7920), .Z(n9090) );
  HS65_LL_NOR3AX2 U15931 ( .A(n8819), .B(n8176), .C(n8804), .Z(n9087) );
  HS65_LL_NOR4ABX2 U15932 ( .A(n8447), .B(n8472), .C(n8775), .D(n8788), .Z(
        n9088) );
  HS65_LL_NOR4ABX2 U15933 ( .A(n9029), .B(n9030), .C(n9031), .D(n9032), .Z(
        n7626) );
  HS65_LL_OAI222X2 U15934 ( .A(n7623), .B(n7821), .C(n7619), .D(n8397), .E(
        n7624), .F(n7822), .Z(n9032) );
  HS65_LL_NOR3AX2 U15935 ( .A(n8729), .B(n8153), .C(n8714), .Z(n9029) );
  HS65_LL_NOR4ABX2 U15936 ( .A(n8395), .B(n8420), .C(n8685), .D(n8698), .Z(
        n9030) );
  HS65_LL_NOR2X6 U15937 ( .A(n8254), .B(n8649), .Z(n8076) );
  HS65_LL_NOR2X6 U15938 ( .A(n3112), .B(n3491), .Z(n3507) );
  HS65_LL_NOR2X6 U15939 ( .A(n7675), .B(n7623), .Z(n8728) );
  HS65_LL_NOR2X6 U15940 ( .A(n7713), .B(n7663), .Z(n8818) );
  HS65_LL_CBI4I1X5 U15941 ( .A(n6143), .B(n6070), .C(n6254), .D(n6295), .Z(
        n7247) );
  HS65_LL_CBI4I1X5 U15942 ( .A(n4550), .B(n4477), .C(n4661), .D(n4702), .Z(
        n5655) );
  HS65_LL_NOR2X6 U15943 ( .A(n4685), .B(n4552), .Z(n5057) );
  HS65_LL_NOR2X6 U15944 ( .A(n6278), .B(n6145), .Z(n6650) );
  HS65_LL_NOR2X6 U15945 ( .A(n2860), .B(n2939), .Z(n3443) );
  HS65_LL_NOR2X6 U15946 ( .A(n3183), .B(n3846), .Z(n3843) );
  HS65_LL_NOR2X6 U15947 ( .A(n3252), .B(n3251), .Z(n3276) );
  HS65_LL_NOR2X6 U15948 ( .A(n8155), .B(n7831), .Z(n8409) );
  HS65_LL_NOR2X6 U15949 ( .A(n8178), .B(n7870), .Z(n8461) );
  HS65_LL_NOR2X6 U15950 ( .A(n7623), .B(n8686), .Z(n8411) );
  HS65_LL_NOR2X6 U15951 ( .A(n7663), .B(n8776), .Z(n8463) );
  HS65_LL_NOR2X6 U15952 ( .A(n3615), .B(n3280), .Z(n3260) );
  HS65_LL_NAND2X7 U15953 ( .A(n7861), .B(n7847), .Z(n7963) );
  HS65_LL_NOR2X6 U15954 ( .A(n3033), .B(n3615), .Z(n3616) );
  HS65_LL_NOR2X6 U15955 ( .A(n3198), .B(n2836), .Z(n3862) );
  HS65_LL_NOR2X6 U15956 ( .A(n7992), .B(n7971), .Z(n8091) );
  HS65_LL_NOR2X6 U15957 ( .A(n7947), .B(n8029), .Z(n8574) );
  HS65_LL_NOR2X6 U15958 ( .A(n5028), .B(n4661), .Z(n4719) );
  HS65_LL_NOR2X6 U15959 ( .A(n6621), .B(n6254), .Z(n6312) );
  HS65_LL_NOR2X6 U15960 ( .A(n4460), .B(n5265), .Z(n5318) );
  HS65_LL_NOR2X6 U15961 ( .A(n6053), .B(n6857), .Z(n6910) );
  HS65_LL_NOR2X6 U15962 ( .A(n4525), .B(n5148), .Z(n5202) );
  HS65_LL_NOR2X6 U15963 ( .A(n6118), .B(n6740), .Z(n6794) );
  HS65_LL_NOR2X6 U15964 ( .A(n4661), .B(n4667), .Z(n5112) );
  HS65_LL_NOR2X6 U15965 ( .A(n6254), .B(n6260), .Z(n6705) );
  HS65_LL_CBI4I1X5 U15966 ( .A(n2956), .B(n2859), .C(n3061), .D(n3435), .Z(
        n4056) );
  HS65_LL_AOI12X2 U15967 ( .A(n7749), .B(n8254), .C(n7993), .Z(n8493) );
  HS65_LL_NOR2X6 U15968 ( .A(n4670), .B(n4551), .Z(n4718) );
  HS65_LL_NOR2X6 U15969 ( .A(n6263), .B(n6144), .Z(n6311) );
  HS65_LL_NAND2X7 U15970 ( .A(n1932), .B(n1931), .Z(n1937) );
  HS65_LL_NAND2X7 U15971 ( .A(n7943), .B(n7948), .Z(n8031) );
  HS65_LL_AOI12X2 U15972 ( .A(n4509), .B(n5382), .C(n5380), .Z(n5558) );
  HS65_LL_AOI12X2 U15973 ( .A(n4448), .B(n5267), .C(n5265), .Z(n5536) );
  HS65_LL_AOI12X2 U15974 ( .A(n4809), .B(n5150), .C(n5148), .Z(n5493) );
  HS65_LL_AOI12X2 U15975 ( .A(n6102), .B(n6974), .C(n6972), .Z(n7150) );
  HS65_LL_AOI12X2 U15976 ( .A(n6402), .B(n6742), .C(n6740), .Z(n7085) );
  HS65_LL_AOI12X2 U15977 ( .A(n6041), .B(n6859), .C(n6857), .Z(n7128) );
  HS65_LL_NOR2X6 U15978 ( .A(n7657), .B(n8173), .Z(n7877) );
  HS65_LL_NOR2X6 U15979 ( .A(n7636), .B(n8150), .Z(n7838) );
  HS65_LL_NAND2X7 U15980 ( .A(n2837), .B(n2992), .Z(n2834) );
  HS65_LL_NAND2X7 U15981 ( .A(n2889), .B(n2981), .Z(n2886) );
  HS65_LL_NAND2X7 U15982 ( .A(n3116), .B(n3464), .Z(n2869) );
  HS65_LL_NOR2X6 U15983 ( .A(n7652), .B(n7656), .Z(n8793) );
  HS65_LL_NOR2X6 U15984 ( .A(n7632), .B(n7619), .Z(n8703) );
  HS65_LL_NOR2X6 U15985 ( .A(n3450), .B(n3114), .Z(n3463) );
  HS65_LL_NAND2X7 U15986 ( .A(n2308), .B(n2307), .Z(n2313) );
  HS65_LL_NOR2X6 U15987 ( .A(n3116), .B(n2957), .Z(n3512) );
  HS65_LL_NOR2X6 U15988 ( .A(n3069), .B(n2859), .Z(n3102) );
  HS65_LL_NOR2X6 U15989 ( .A(n2838), .B(n2997), .Z(n3385) );
  HS65_LL_NOR2X6 U15990 ( .A(n3158), .B(n3299), .Z(n3156) );
  HS65_LL_NOR2X6 U15991 ( .A(n3225), .B(n3251), .Z(n3028) );
  HS65_LL_NOR2X6 U15992 ( .A(n8034), .B(n8357), .Z(n8583) );
  HS65_LL_NAND4ABX3 U15993 ( .A(n6418), .B(n6419), .C(n6420), .D(n6421), .Z(
        n6214) );
  HS65_LL_NAND4ABX3 U15994 ( .A(n6449), .B(n6450), .C(n6451), .D(n6452), .Z(
        n6419) );
  HS65_LL_NOR4ABX2 U15995 ( .A(n6422), .B(n6423), .C(n6424), .D(n6425), .Z(
        n6421) );
  HS65_LL_MX41X7 U15996 ( .D0(n6114), .S0(n515), .D1(n490), .S1(n521), .D2(
        n523), .S2(n498), .D3(n502), .S3(n518), .Z(n6418) );
  HS65_LL_NAND4ABX3 U15997 ( .A(n4825), .B(n4826), .C(n4827), .D(n4828), .Z(
        n4621) );
  HS65_LL_NAND4ABX3 U15998 ( .A(n4856), .B(n4857), .C(n4858), .D(n4859), .Z(
        n4826) );
  HS65_LL_NOR4ABX2 U15999 ( .A(n4829), .B(n4830), .C(n4831), .D(n4832), .Z(
        n4828) );
  HS65_LL_MX41X7 U16000 ( .D0(n4521), .S0(n691), .D1(n666), .S1(n697), .D2(
        n699), .S2(n674), .D3(n678), .S3(n694), .Z(n4825) );
  HS65_LL_OAI21X3 U16001 ( .A(n3450), .B(n3060), .C(n4049), .Z(n4048) );
  HS65_LL_OAI21X3 U16002 ( .A(n190), .B(n192), .C(n209), .Z(n4049) );
  HS65_LL_NAND2X7 U16003 ( .A(n1556), .B(n1555), .Z(n1561) );
  HS65_LL_NAND4ABX3 U16004 ( .A(n8327), .B(n8328), .C(n8329), .D(n8330), .Z(
        n7939) );
  HS65_LL_OAI222X2 U16005 ( .A(n8339), .B(n7948), .C(n8049), .D(n8057), .E(
        n7767), .F(n7769), .Z(n8328) );
  HS65_LL_NOR4ABX2 U16006 ( .A(n8331), .B(n8332), .C(n8333), .D(n8334), .Z(
        n8330) );
  HS65_LL_NAND3X5 U16007 ( .A(n8340), .B(n8341), .C(n8342), .Z(n8327) );
  HS65_LL_NOR2X6 U16008 ( .A(n6402), .B(n6221), .Z(n6449) );
  HS65_LL_NOR2X6 U16009 ( .A(n4809), .B(n4628), .Z(n4856) );
  HS65_LL_NAND2X7 U16010 ( .A(n2958), .B(n2957), .Z(n2963) );
  HS65_LL_NAND2X7 U16011 ( .A(n3185), .B(n3183), .Z(n3190) );
  HS65_LL_NOR2X6 U16012 ( .A(n7632), .B(n8145), .Z(n8749) );
  HS65_LL_NOR2X6 U16013 ( .A(n7652), .B(n8168), .Z(n8839) );
  HS65_LL_NOR2X6 U16014 ( .A(n4448), .B(n4747), .Z(n4920) );
  HS65_LL_NOR2X6 U16015 ( .A(n4509), .B(n4773), .Z(n4973) );
  HS65_LL_NOR2X6 U16016 ( .A(n4809), .B(n4627), .Z(n4845) );
  HS65_LL_NOR2X6 U16017 ( .A(n6102), .B(n6366), .Z(n6566) );
  HS65_LL_NOR2X6 U16018 ( .A(n6402), .B(n6220), .Z(n6438) );
  HS65_LL_NOR2X6 U16019 ( .A(n6041), .B(n6327), .Z(n6513) );
  HS65_LL_IVX9 U16020 ( .A(n3061), .Z(n224) );
  HS65_LL_NOR2X6 U16021 ( .A(n7905), .B(n8173), .Z(n7876) );
  HS65_LL_NOR2X6 U16022 ( .A(n7807), .B(n8150), .Z(n7837) );
  HS65_LL_NOR2X6 U16023 ( .A(n2890), .B(n2968), .Z(n3327) );
  HS65_LL_NOR2X6 U16024 ( .A(n2838), .B(n2993), .Z(n3381) );
  HS65_LL_NOR2X6 U16025 ( .A(n7664), .B(n7714), .Z(n8805) );
  HS65_LL_NOR2X6 U16026 ( .A(n7624), .B(n7676), .Z(n8715) );
  HS65_LL_IVX9 U16027 ( .A(n2914), .Z(n153) );
  HS65_LL_OAI21X3 U16028 ( .A(n2940), .B(n3069), .C(n3070), .Z(n3068) );
  HS65_LL_IVX9 U16029 ( .A(n6302), .Z(n556) );
  HS65_LL_IVX9 U16030 ( .A(n4709), .Z(n34) );
  HS65_LL_NOR2X6 U16031 ( .A(n3115), .B(n3067), .Z(n3444) );
  HS65_LL_NAND2X7 U16032 ( .A(n4500), .B(n4610), .Z(n4497) );
  HS65_LL_NAND2X7 U16033 ( .A(n4461), .B(n4593), .Z(n4458) );
  HS65_LL_NAND2X7 U16034 ( .A(n6093), .B(n6203), .Z(n6090) );
  HS65_LL_NAND2X7 U16035 ( .A(n5496), .B(n5135), .Z(n4527) );
  HS65_LL_NAND2X7 U16036 ( .A(n7088), .B(n6727), .Z(n6120) );
  HS65_LL_NAND2X7 U16037 ( .A(n6054), .B(n6186), .Z(n6051) );
  HS65_LL_NAND2X7 U16038 ( .A(n5502), .B(n5472), .Z(n5077) );
  HS65_LL_NAND2X7 U16039 ( .A(n7094), .B(n7064), .Z(n6670) );
  HS65_LL_NOR2X6 U16040 ( .A(n6441), .B(n6442), .Z(n6411) );
  HS65_LL_NOR2X6 U16041 ( .A(n4848), .B(n4849), .Z(n4818) );
  HS65_LL_IVX9 U16042 ( .A(n7632), .Z(n584) );
  HS65_LL_IVX9 U16043 ( .A(n7652), .Z(n104) );
  HS65_LL_NOR2X6 U16044 ( .A(n3326), .B(n3141), .Z(n3310) );
  HS65_LL_NAND2X7 U16045 ( .A(n3158), .B(n3157), .Z(n3163) );
  HS65_LL_NOR2X6 U16046 ( .A(n6441), .B(n6126), .Z(n6764) );
  HS65_LL_NOR2X6 U16047 ( .A(n4848), .B(n4533), .Z(n5172) );
  HS65_LL_NOR2X6 U16048 ( .A(n4456), .B(n4586), .Z(n5288) );
  HS65_LL_NOR2X6 U16049 ( .A(n4495), .B(n4603), .Z(n5403) );
  HS65_LL_NOR2X6 U16050 ( .A(n6049), .B(n6179), .Z(n6880) );
  HS65_LL_NOR2X6 U16051 ( .A(n6088), .B(n6196), .Z(n6995) );
  HS65_LL_NOR2X6 U16052 ( .A(n6302), .B(n6304), .Z(n6271) );
  HS65_LL_NOR2X6 U16053 ( .A(n4709), .B(n4711), .Z(n4678) );
  HS65_LL_NAND2X7 U16054 ( .A(n3271), .B(n3588), .Z(n2912) );
  HS65_LL_NAND4ABX3 U16055 ( .A(n5830), .B(n5831), .C(n5832), .D(n5833), .Z(
        n4451) );
  HS65_LL_OAI222X2 U16056 ( .A(n4460), .B(n4876), .C(n5267), .D(n4883), .E(
        n4453), .F(n4593), .Z(n5830) );
  HS65_LL_NOR3AX2 U16057 ( .A(n5244), .B(n5262), .C(n5306), .Z(n5833) );
  HS65_LL_NAND4ABX3 U16058 ( .A(n4760), .B(n4920), .C(n5347), .D(n5280), .Z(
        n5831) );
  HS65_LL_NAND4ABX3 U16059 ( .A(n5889), .B(n5890), .C(n5891), .D(n5892), .Z(
        n4512) );
  HS65_LL_OAI222X2 U16060 ( .A(n4499), .B(n4988), .C(n5382), .D(n4995), .E(
        n4492), .F(n4610), .Z(n5889) );
  HS65_LL_NOR3AX2 U16061 ( .A(n5359), .B(n5377), .C(n5421), .Z(n5892) );
  HS65_LL_NAND4ABX3 U16062 ( .A(n4787), .B(n4973), .C(n5462), .D(n5395), .Z(
        n5890) );
  HS65_LL_NAND4ABX3 U16063 ( .A(n5774), .B(n5775), .C(n5776), .D(n5777), .Z(
        n5675) );
  HS65_LL_OAI222X2 U16064 ( .A(n4525), .B(n4862), .C(n5150), .D(n4869), .E(
        n4850), .F(n5135), .Z(n5774) );
  HS65_LL_NOR3AX2 U16065 ( .A(n5126), .B(n5145), .C(n5190), .Z(n5777) );
  HS65_LL_NAND4ABX3 U16066 ( .A(n4641), .B(n4845), .C(n5232), .D(n5163), .Z(
        n5775) );
  HS65_LL_NAND4ABX3 U16067 ( .A(n7481), .B(n7482), .C(n7483), .D(n7484), .Z(
        n6105) );
  HS65_LL_OAI222X2 U16068 ( .A(n6092), .B(n6581), .C(n6974), .D(n6588), .E(
        n6085), .F(n6203), .Z(n7481) );
  HS65_LL_NOR3AX2 U16069 ( .A(n6951), .B(n6969), .C(n7013), .Z(n7484) );
  HS65_LL_NAND4ABX3 U16070 ( .A(n6380), .B(n6566), .C(n7054), .D(n6987), .Z(
        n7482) );
  HS65_LL_NAND4ABX3 U16071 ( .A(n7366), .B(n7367), .C(n7368), .D(n7369), .Z(
        n7267) );
  HS65_LL_OAI222X2 U16072 ( .A(n6118), .B(n6455), .C(n6742), .D(n6462), .E(
        n6443), .F(n6727), .Z(n7366) );
  HS65_LL_NOR3AX2 U16073 ( .A(n6718), .B(n6737), .C(n6782), .Z(n7369) );
  HS65_LL_NAND4ABX3 U16074 ( .A(n6234), .B(n6438), .C(n6824), .D(n6755), .Z(
        n7367) );
  HS65_LL_NAND4ABX3 U16075 ( .A(n7422), .B(n7423), .C(n7424), .D(n7425), .Z(
        n6044) );
  HS65_LL_OAI222X2 U16076 ( .A(n6053), .B(n6469), .C(n6859), .D(n6476), .E(
        n6046), .F(n6186), .Z(n7422) );
  HS65_LL_NOR3AX2 U16077 ( .A(n6836), .B(n6854), .C(n6898), .Z(n7425) );
  HS65_LL_NAND4ABX3 U16078 ( .A(n6341), .B(n6513), .C(n6939), .D(n6872), .Z(
        n7423) );
  HS65_LL_CBI4I1X5 U16079 ( .A(n4626), .B(n4533), .C(n4862), .D(n4840), .Z(
        n5685) );
  HS65_LL_CBI4I1X5 U16080 ( .A(n6219), .B(n6126), .C(n6455), .D(n6433), .Z(
        n7277) );
  HS65_LL_NAND4ABX3 U16081 ( .A(n2945), .B(n2946), .C(n2947), .D(n2948), .Z(
        n2866) );
  HS65_LL_NOR3AX2 U16082 ( .A(n2953), .B(n2954), .C(n2955), .Z(n2947) );
  HS65_LL_NOR4ABX2 U16083 ( .A(n2949), .B(n2950), .C(n2951), .D(n2952), .Z(
        n2948) );
  HS65_LL_OAI212X5 U16084 ( .A(n2956), .B(n2957), .C(n2932), .D(n2958), .E(
        n2959), .Z(n2946) );
  HS65_LL_NAND4ABX3 U16085 ( .A(n3172), .B(n3173), .C(n3174), .D(n3175), .Z(
        n2989) );
  HS65_LL_NOR4ABX2 U16086 ( .A(n3176), .B(n3177), .C(n3178), .D(n3179), .Z(
        n3175) );
  HS65_LL_NOR3AX2 U16087 ( .A(n3180), .B(n3181), .C(n3182), .Z(n3174) );
  HS65_LL_OAI212X5 U16088 ( .A(n2832), .B(n3183), .C(n3184), .D(n3185), .E(
        n3186), .Z(n3173) );
  HS65_LL_NAND4ABX3 U16089 ( .A(n3146), .B(n3147), .C(n3148), .D(n3149), .Z(
        n2978) );
  HS65_LL_NOR3AX2 U16090 ( .A(n3154), .B(n3155), .C(n3156), .Z(n3148) );
  HS65_LL_NOR4ABX2 U16091 ( .A(n3150), .B(n3151), .C(n3152), .D(n3153), .Z(
        n3149) );
  HS65_LL_OAI212X5 U16092 ( .A(n2884), .B(n3157), .C(n3134), .D(n3158), .E(
        n3159), .Z(n3147) );
  HS65_LL_NAND4ABX3 U16093 ( .A(n8377), .B(n8378), .C(n8379), .D(n8380), .Z(
        n8140) );
  HS65_LL_NAND4ABX3 U16094 ( .A(n7788), .B(n8401), .C(n8402), .D(n8403), .Z(
        n8378) );
  HS65_LL_MX41X7 U16095 ( .D0(n606), .S0(n7699), .D1(n583), .S1(n612), .D2(
        n599), .S2(n592), .D3(n586), .S3(n609), .Z(n8377) );
  HS65_LL_NOR4ABX2 U16096 ( .A(n8381), .B(n8382), .C(n8383), .D(n8384), .Z(
        n8380) );
  HS65_LL_NAND4ABX3 U16097 ( .A(n8429), .B(n8430), .C(n8431), .D(n8432), .Z(
        n8163) );
  HS65_LL_NAND4ABX3 U16098 ( .A(n7887), .B(n8453), .C(n8454), .D(n8455), .Z(
        n8430) );
  HS65_LL_MX41X7 U16099 ( .D0(n126), .S0(n7737), .D1(n103), .S1(n132), .D2(
        n119), .S2(n112), .D3(n106), .S3(n129), .Z(n8429) );
  HS65_LL_NOR4ABX2 U16100 ( .A(n8433), .B(n8434), .C(n8435), .D(n8436), .Z(
        n8432) );
  HS65_LL_NOR2X6 U16101 ( .A(n4988), .B(n4994), .Z(n4503) );
  HS65_LL_NOR2X6 U16102 ( .A(n4876), .B(n4882), .Z(n4464) );
  HS65_LL_NOR2X6 U16103 ( .A(n6581), .B(n6587), .Z(n6096) );
  HS65_LL_NOR2X6 U16104 ( .A(n4862), .B(n4868), .Z(n5218) );
  HS65_LL_NOR2X6 U16105 ( .A(n6455), .B(n6461), .Z(n6810) );
  HS65_LL_NOR2X6 U16106 ( .A(n6469), .B(n6475), .Z(n6057) );
  HS65_LL_NOR2X6 U16107 ( .A(n3982), .B(n3047), .Z(n3612) );
  HS65_LL_NAND2X7 U16108 ( .A(n44), .B(n4481), .Z(n5046) );
  HS65_LL_NAND2X7 U16109 ( .A(n566), .B(n6074), .Z(n6639) );
  HS65_LL_NOR2X6 U16110 ( .A(n8254), .B(n8106), .Z(n8101) );
  HS65_LL_NAND2X7 U16111 ( .A(n119), .B(n7737), .Z(n8790) );
  HS65_LL_NOR2X6 U16112 ( .A(n2957), .B(n3491), .Z(n3487) );
  HS65_LL_IVX9 U16113 ( .A(n3225), .Z(n145) );
  HS65_LL_AOI12X2 U16114 ( .A(n7836), .B(n8005), .C(n7632), .Z(n8004) );
  HS65_LL_AOI12X2 U16115 ( .A(n7875), .B(n8018), .C(n7652), .Z(n8017) );
  HS65_LL_NOR2X6 U16116 ( .A(n4775), .B(n4508), .Z(n5410) );
  HS65_LL_NOR2X6 U16117 ( .A(n4629), .B(n4654), .Z(n5179) );
  HS65_LL_NOR2X6 U16118 ( .A(n6222), .B(n6247), .Z(n6771) );
  HS65_LL_NOR2X6 U16119 ( .A(n6368), .B(n6101), .Z(n7002) );
  HS65_LL_NAND2X7 U16120 ( .A(n132), .B(n7737), .Z(n7890) );
  HS65_LL_NAND2X7 U16121 ( .A(n8049), .B(n8048), .Z(n7761) );
  HS65_LL_NOR2X6 U16122 ( .A(n3225), .B(n3984), .Z(n3553) );
  HS65_LL_NOR2X6 U16123 ( .A(n3615), .B(n3984), .Z(n3277) );
  HS65_LL_NOR2X6 U16124 ( .A(n5267), .B(n5532), .Z(n5263) );
  HS65_LL_NOR2X6 U16125 ( .A(n5382), .B(n5554), .Z(n5378) );
  HS65_LL_NOR2X6 U16126 ( .A(n5150), .B(n5579), .Z(n5146) );
  HS65_LL_NOR2X6 U16127 ( .A(n6859), .B(n7124), .Z(n6855) );
  HS65_LL_NOR2X6 U16128 ( .A(n6974), .B(n7146), .Z(n6970) );
  HS65_LL_NOR2X6 U16129 ( .A(n6742), .B(n7171), .Z(n6738) );
  HS65_LL_CBI4I1X5 U16130 ( .A(n2832), .B(n2997), .C(n3406), .D(n3793), .Z(
        n4295) );
  HS65_LL_IVX9 U16131 ( .A(n4809), .Z(n668) );
  HS65_LL_IVX9 U16132 ( .A(n6402), .Z(n492) );
  HS65_LL_NOR2X6 U16133 ( .A(n4922), .B(n5604), .Z(n4736) );
  HS65_LL_NOR2X6 U16134 ( .A(n4975), .B(n5629), .Z(n4797) );
  HS65_LL_NOR2X6 U16135 ( .A(n6568), .B(n7221), .Z(n6390) );
  HS65_LL_NOR2X6 U16136 ( .A(n6515), .B(n7196), .Z(n6351) );
  HS65_LL_NOR2X6 U16137 ( .A(n6440), .B(n7170), .Z(n6244) );
  HS65_LL_NOR2X6 U16138 ( .A(n4847), .B(n5578), .Z(n4651) );
  HS65_LL_CBI4I1X5 U16139 ( .A(n3406), .B(n3185), .C(n2836), .D(n3831), .Z(
        n3830) );
  HS65_LL_NOR2X6 U16140 ( .A(n5026), .B(n4711), .Z(n4554) );
  HS65_LL_NOR2X6 U16141 ( .A(n6619), .B(n6304), .Z(n6147) );
  HS65_LL_NAND2X7 U16142 ( .A(n7981), .B(n7980), .Z(n7743) );
  HS65_LL_NOR2X6 U16143 ( .A(n6278), .B(n7094), .Z(n6148) );
  HS65_LL_NOR2X6 U16144 ( .A(n4685), .B(n5502), .Z(n4555) );
  HS65_LL_AOI12X2 U16145 ( .A(n1881), .B(n2071), .C(n2069), .Z(n2145) );
  HS65_LL_AOI12X2 U16146 ( .A(n1129), .B(n1319), .C(n1317), .Z(n1393) );
  HS65_LL_AOI12X2 U16147 ( .A(n2875), .B(n3731), .C(n3343), .Z(n3951) );
  HS65_LL_AOI12X2 U16148 ( .A(n6116), .B(n6117), .C(n6118), .Z(n6115) );
  HS65_LL_AOI12X2 U16149 ( .A(n4523), .B(n4524), .C(n4525), .Z(n4522) );
  HS65_LL_AOI12X2 U16150 ( .A(n4462), .B(n4591), .C(n4460), .Z(n4590) );
  HS65_LL_AOI12X2 U16151 ( .A(n6094), .B(n6201), .C(n6092), .Z(n6200) );
  HS65_LL_AOI12X2 U16152 ( .A(n6055), .B(n6184), .C(n6053), .Z(n6183) );
  HS65_LL_AOI12X2 U16153 ( .A(n4501), .B(n4608), .C(n4499), .Z(n4607) );
  HS65_LL_NAND2X7 U16154 ( .A(n472), .B(n4606), .Z(n5400) );
  HS65_LL_NAND2X7 U16155 ( .A(n255), .B(n4589), .Z(n5285) );
  HS65_LL_NAND2X7 U16156 ( .A(n699), .B(n4521), .Z(n5168) );
  HS65_LL_NAND2X7 U16157 ( .A(n297), .B(n6199), .Z(n6992) );
  HS65_LL_NAND2X7 U16158 ( .A(n523), .B(n6114), .Z(n6760) );
  HS65_LL_AOI12X2 U16159 ( .A(n2257), .B(n2447), .C(n2445), .Z(n2521) );
  HS65_LL_CBI4I1X5 U16160 ( .A(n2276), .B(n2238), .C(n2277), .D(n2278), .Z(
        n2261) );
  HS65_LL_CBI4I1X5 U16161 ( .A(n1900), .B(n1862), .C(n1901), .D(n1902), .Z(
        n1885) );
  HS65_LL_NOR2X6 U16162 ( .A(n4710), .B(n5514), .Z(n4574) );
  HS65_LL_NOR2X6 U16163 ( .A(n6303), .B(n7106), .Z(n6167) );
  HS65_LL_NAND2X7 U16164 ( .A(n2245), .B(n2271), .Z(n2242) );
  HS65_LL_NAND2X7 U16165 ( .A(n1493), .B(n1519), .Z(n1490) );
  HS65_LL_NAND2X7 U16166 ( .A(n1117), .B(n1143), .Z(n1114) );
  HS65_LL_NAND2X7 U16167 ( .A(n1869), .B(n1895), .Z(n1866) );
  HS65_LL_NOR2X6 U16168 ( .A(n4790), .B(n4994), .Z(n4502) );
  HS65_LL_NOR2X6 U16169 ( .A(n4728), .B(n4882), .Z(n4463) );
  HS65_LL_NOR2X6 U16170 ( .A(n6383), .B(n6587), .Z(n6095) );
  HS65_LL_NOR2X6 U16171 ( .A(n4644), .B(n4868), .Z(n5170) );
  HS65_LL_NOR2X6 U16172 ( .A(n6237), .B(n6461), .Z(n6762) );
  HS65_LL_NOR2X6 U16173 ( .A(n6344), .B(n6475), .Z(n6056) );
  HS65_LL_AOI12X2 U16174 ( .A(n1505), .B(n1695), .C(n1693), .Z(n1769) );
  HS65_LL_IVX9 U16175 ( .A(n3406), .Z(n433) );
  HS65_LL_IVX9 U16176 ( .A(n3396), .Z(n415) );
  HS65_LL_IVX9 U16177 ( .A(n3114), .Z(n192) );
  HS65_LL_NOR2X6 U16178 ( .A(n7947), .B(n7942), .Z(n8576) );
  HS65_LL_AOI12X2 U16179 ( .A(n2940), .B(n3491), .C(n3115), .Z(n3898) );
  HS65_LL_IVX9 U16180 ( .A(n6118), .Z(n489) );
  HS65_LL_IVX9 U16181 ( .A(n4525), .Z(n665) );
  HS65_LL_NOR3X4 U16182 ( .A(n4087), .B(n4088), .C(n3906), .Z(n4084) );
  HS65_LL_OAI21X3 U16183 ( .A(n3047), .B(n3034), .C(n4095), .Z(n4087) );
  HS65_LL_NOR2X6 U16184 ( .A(n3042), .B(n3251), .Z(n3645) );
  HS65_LL_NAND2X7 U16185 ( .A(n7874), .B(n7919), .Z(n7872) );
  HS65_LL_NAND2X7 U16186 ( .A(n7835), .B(n7821), .Z(n7833) );
  HS65_LL_NOR2X6 U16187 ( .A(n7851), .B(n7971), .Z(n8306) );
  HS65_LL_IVX9 U16188 ( .A(n7870), .Z(n124) );
  HS65_LL_NOR2X6 U16189 ( .A(n3033), .B(n2917), .Z(n3555) );
  HS65_LL_IVX9 U16190 ( .A(n6441), .Z(n513) );
  HS65_LL_IVX9 U16191 ( .A(n4848), .Z(n689) );
  HS65_LL_IVX9 U16192 ( .A(n6462), .Z(n509) );
  HS65_LL_IVX9 U16193 ( .A(n4883), .Z(n259) );
  HS65_LL_IVX9 U16194 ( .A(n4869), .Z(n685) );
  HS65_LL_NAND3X5 U16195 ( .A(n6254), .B(n7093), .C(n6158), .Z(n7108) );
  HS65_LL_NAND3X5 U16196 ( .A(n4661), .B(n5501), .C(n4565), .Z(n5516) );
  HS65_LL_OAI21X3 U16197 ( .A(n5508), .B(n4660), .C(n5643), .Z(n5642) );
  HS65_LL_OAI21X3 U16198 ( .A(n11), .B(n14), .C(n39), .Z(n5643) );
  HS65_LL_OAI21X3 U16199 ( .A(n7100), .B(n6253), .C(n7235), .Z(n7234) );
  HS65_LL_OAI21X3 U16200 ( .A(n533), .B(n536), .C(n561), .Z(n7235) );
  HS65_LL_OAI21X3 U16201 ( .A(n7767), .B(n8313), .C(n8314), .Z(n8312) );
  HS65_LL_IVX9 U16202 ( .A(n3251), .Z(n167) );
  HS65_LL_NAND2X7 U16203 ( .A(n4748), .B(n4747), .Z(n4757) );
  HS65_LL_NAND2X7 U16204 ( .A(n4774), .B(n4773), .Z(n4784) );
  HS65_LL_NAND2X7 U16205 ( .A(n4628), .B(n4627), .Z(n4638) );
  HS65_LL_NAND2X7 U16206 ( .A(n6328), .B(n6327), .Z(n6338) );
  HS65_LL_NAND2X7 U16207 ( .A(n6367), .B(n6366), .Z(n6377) );
  HS65_LL_NAND2X7 U16208 ( .A(n6221), .B(n6220), .Z(n6231) );
  HS65_LL_IVX9 U16209 ( .A(n2915), .Z(n164) );
  HS65_LL_CBI4I1X5 U16210 ( .A(n8363), .B(n8049), .C(n8540), .D(n8541), .Z(
        n8539) );
  HS65_LL_NOR2X6 U16211 ( .A(n7768), .B(n8039), .Z(n8610) );
  HS65_LL_NOR4ABX2 U16212 ( .A(n3263), .B(n3264), .C(n3265), .D(n3266), .Z(
        n2906) );
  HS65_LL_OAI222X2 U16213 ( .A(n3269), .B(n3270), .C(n3271), .D(n3253), .E(
        n3047), .F(n3043), .Z(n3265) );
  HS65_LL_OAI212X5 U16214 ( .A(n3267), .B(n3054), .C(n3224), .D(n3042), .E(
        n3268), .Z(n3266) );
  HS65_LL_NOR3AX2 U16215 ( .A(n3272), .B(n3273), .C(n3274), .Z(n3264) );
  HS65_LL_NOR2X6 U16216 ( .A(n3157), .B(n3299), .Z(n3727) );
  HS65_LL_NOR2X6 U16217 ( .A(n2890), .B(n2972), .Z(n3331) );
  HS65_LL_NOR4ABX2 U16218 ( .A(n3390), .B(n3391), .C(n3392), .D(n3393), .Z(
        n2986) );
  HS65_LL_OAI222X2 U16219 ( .A(n3396), .B(n3397), .C(n2837), .D(n2829), .E(
        n3197), .F(n3193), .Z(n3392) );
  HS65_LL_NOR3X4 U16220 ( .A(n3398), .B(n3399), .C(n3400), .Z(n3391) );
  HS65_LL_OAI212X5 U16221 ( .A(n3394), .B(n2846), .C(n3192), .D(n2838), .E(
        n3395), .Z(n3393) );
  HS65_LL_NOR4ABX2 U16222 ( .A(n3107), .B(n3108), .C(n3109), .D(n3110), .Z(
        n2863) );
  HS65_LL_OAI222X2 U16223 ( .A(n3114), .B(n3115), .C(n3116), .D(n3097), .E(
        n2931), .F(n2927), .Z(n3109) );
  HS65_LL_NOR3X4 U16224 ( .A(n3117), .B(n3118), .C(n3119), .Z(n3108) );
  HS65_LL_OAI212X5 U16225 ( .A(n3111), .B(n3112), .C(n2926), .D(n3069), .E(
        n3113), .Z(n3110) );
  HS65_LL_NOR2X6 U16226 ( .A(n6621), .B(n6144), .Z(n6156) );
  HS65_LL_NOR2X6 U16227 ( .A(n5028), .B(n4551), .Z(n4563) );
  HS65_LL_NOR2X6 U16228 ( .A(n5382), .B(n4495), .Z(n4981) );
  HS65_LL_NOR2X6 U16229 ( .A(n5267), .B(n4456), .Z(n4928) );
  HS65_LL_NOR2X6 U16230 ( .A(n6974), .B(n6088), .Z(n6574) );
  HS65_LL_NOR2X6 U16231 ( .A(n5150), .B(n4848), .Z(n4855) );
  HS65_LL_NOR2X6 U16232 ( .A(n6742), .B(n6441), .Z(n6448) );
  HS65_LL_NOR2X6 U16233 ( .A(n6859), .B(n6049), .Z(n6521) );
  HS65_LL_NOR4ABX2 U16234 ( .A(n8349), .B(n8350), .C(n8351), .D(n8352), .Z(
        n7936) );
  HS65_LL_OAI212X5 U16235 ( .A(n8356), .B(n8357), .C(n8028), .D(n8313), .E(
        n8358), .Z(n8351) );
  HS65_LL_AOI222X2 U16236 ( .A(n333), .B(n352), .C(n342), .D(n332), .E(n335), 
        .F(n347), .Z(n8349) );
  HS65_LL_NAND3AX6 U16237 ( .A(n8353), .B(n8354), .C(n8355), .Z(n8352) );
  HS65_LL_NOR2X6 U16238 ( .A(n4551), .B(n4667), .Z(n4564) );
  HS65_LL_NOR2X6 U16239 ( .A(n6144), .B(n6260), .Z(n6157) );
  HS65_LL_NOR2X6 U16240 ( .A(n2957), .B(n2856), .Z(n3442) );
  HS65_LL_IVX9 U16241 ( .A(n7660), .Z(n99) );
  HS65_LL_IVX9 U16242 ( .A(n7620), .Z(n579) );
  HS65_LL_NOR2X6 U16243 ( .A(n3615), .B(n3251), .Z(n3254) );
  HS65_LL_IVX9 U16244 ( .A(n4627), .Z(n692) );
  HS65_LL_IVX9 U16245 ( .A(n6220), .Z(n516) );
  HS65_LL_NAND2X7 U16246 ( .A(n3491), .B(n2856), .Z(n3417) );
  HS65_LL_CBI4I1X5 U16247 ( .A(n1693), .B(n1485), .C(n1537), .D(n1796), .Z(
        n1774) );
  HS65_LL_AO12X9 U16248 ( .A(n1544), .B(n1525), .C(n1745), .Z(n1796) );
  HS65_LL_NOR2X6 U16249 ( .A(n4567), .B(n4711), .Z(n5088) );
  HS65_LL_NOR2X6 U16250 ( .A(n6160), .B(n6304), .Z(n6681) );
  HS65_LL_NOR2X6 U16251 ( .A(n3269), .B(n3286), .Z(n3568) );
  HS65_LL_NOR2X6 U16252 ( .A(n7870), .B(n8776), .Z(n8452) );
  HS65_LL_NOR2X6 U16253 ( .A(n7831), .B(n8686), .Z(n8400) );
  HS65_LL_NOR2X6 U16254 ( .A(n5028), .B(n4709), .Z(n4717) );
  HS65_LL_NOR2X6 U16255 ( .A(n6621), .B(n6302), .Z(n6310) );
  HS65_LL_NOR2X6 U16256 ( .A(n8397), .B(n7623), .Z(n8134) );
  HS65_LL_IVX9 U16257 ( .A(n8145), .Z(n605) );
  HS65_LL_IVX9 U16258 ( .A(n8168), .Z(n125) );
  HS65_LL_IVX9 U16259 ( .A(n5501), .Z(n47) );
  HS65_LL_IVX9 U16260 ( .A(n7093), .Z(n569) );
  HS65_LL_NOR4ABX2 U16261 ( .A(n7976), .B(n7977), .C(n7978), .D(n7979), .Z(
        n7855) );
  HS65_LL_NAND4ABX3 U16262 ( .A(n7983), .B(n7984), .C(n7985), .D(n7986), .Z(
        n7978) );
  HS65_LL_NOR3X4 U16263 ( .A(n7747), .B(n7990), .C(n7991), .Z(n7976) );
  HS65_LL_OAI212X5 U16264 ( .A(n7980), .B(n7861), .C(n7981), .D(n7966), .E(
        n7982), .Z(n7979) );
  HS65_LL_NOR4ABX2 U16265 ( .A(n8044), .B(n8045), .C(n8046), .D(n8047), .Z(
        n7937) );
  HS65_LL_NOR3X4 U16266 ( .A(n8059), .B(n8060), .C(n8061), .Z(n8044) );
  HS65_LL_OAI212X5 U16267 ( .A(n8048), .B(n7943), .C(n8049), .D(n8034), .E(
        n8050), .Z(n8047) );
  HS65_LL_NAND4ABX3 U16268 ( .A(n8051), .B(n8052), .C(n8053), .D(n8054), .Z(
        n8046) );
  HS65_LL_NOR2X6 U16269 ( .A(n7713), .B(n7905), .Z(n8792) );
  HS65_LL_NOR2X6 U16270 ( .A(n7675), .B(n7807), .Z(n8702) );
  HS65_LL_AOI12X2 U16271 ( .A(n2845), .B(n3846), .C(n3397), .Z(n3971) );
  HS65_LL_IVX9 U16272 ( .A(n5026), .Z(n36) );
  HS65_LL_IVX9 U16273 ( .A(n6619), .Z(n558) );
  HS65_LL_NOR2X6 U16274 ( .A(n7947), .B(n8630), .Z(n8558) );
  HS65_LL_NOR2X6 U16275 ( .A(n7846), .B(n8649), .Z(n8256) );
  HS65_LL_NAND2X7 U16276 ( .A(n8556), .B(n7948), .Z(n8498) );
  HS65_LL_NOR2X6 U16277 ( .A(n5382), .B(n4508), .Z(n5402) );
  HS65_LL_NOR2X6 U16278 ( .A(n6974), .B(n6101), .Z(n6994) );
  HS65_LL_NOR2X6 U16279 ( .A(n5267), .B(n4447), .Z(n5287) );
  HS65_LL_NOR2X6 U16280 ( .A(n6742), .B(n6247), .Z(n6763) );
  HS65_LL_NOR2X6 U16281 ( .A(n5150), .B(n4654), .Z(n5171) );
  HS65_LL_NOR2X6 U16282 ( .A(n3293), .B(n3299), .Z(n2892) );
  HS65_LL_NOR2X6 U16283 ( .A(n7636), .B(n8686), .Z(n8401) );
  HS65_LL_NOR2X6 U16284 ( .A(n7657), .B(n8776), .Z(n8453) );
  HS65_LL_IVX9 U16285 ( .A(n2831), .Z(n439) );
  HS65_LL_NOR4ABX2 U16286 ( .A(n8293), .B(n8294), .C(n8295), .D(n8296), .Z(
        n8069) );
  HS65_LL_NAND4ABX3 U16287 ( .A(n8297), .B(n8298), .C(n8299), .D(n8300), .Z(
        n8296) );
  HS65_LL_NOR3X4 U16288 ( .A(n8305), .B(n8306), .C(n8307), .Z(n8294) );
  HS65_LL_OAI212X5 U16289 ( .A(n8301), .B(n8302), .C(n8303), .D(n7750), .E(
        n8304), .Z(n8295) );
  HS65_LL_NOR2X6 U16290 ( .A(n5028), .B(n5501), .Z(n5024) );
  HS65_LL_NOR2X6 U16291 ( .A(n6621), .B(n7093), .Z(n6617) );
  HS65_LL_IVX9 U16292 ( .A(n2957), .Z(n215) );
  HS65_LL_IVX9 U16293 ( .A(n3183), .Z(n437) );
  HS65_LL_IVX9 U16294 ( .A(n3982), .Z(n180) );
  HS65_LL_IVX9 U16295 ( .A(n3271), .Z(n148) );
  HS65_LL_IVX9 U16296 ( .A(n3984), .Z(n165) );
  HS65_LL_NOR2X6 U16297 ( .A(n3033), .B(n3053), .Z(n3581) );
  HS65_LL_NOR2X6 U16298 ( .A(n3033), .B(n2914), .Z(n3569) );
  HS65_LL_OAI21X3 U16299 ( .A(n7749), .B(n8067), .C(n8068), .Z(n8066) );
  HS65_LL_NAND3X5 U16300 ( .A(n3982), .B(n3280), .C(n3041), .Z(n3995) );
  HS65_LL_NOR2X6 U16301 ( .A(n8369), .B(n8049), .Z(n8061) );
  HS65_LL_NAND4ABX3 U16302 ( .A(n8094), .B(n8095), .C(n8096), .D(n8097), .Z(
        n7857) );
  HS65_LL_OAI222X2 U16303 ( .A(n8106), .B(n7847), .C(n7981), .D(n7992), .E(
        n7749), .F(n7751), .Z(n8095) );
  HS65_LL_NOR4ABX2 U16304 ( .A(n8098), .B(n8099), .C(n8100), .D(n8101), .Z(
        n8097) );
  HS65_LL_NAND3X5 U16305 ( .A(n8107), .B(n8108), .C(n8109), .Z(n8094) );
  HS65_LL_NOR2X6 U16306 ( .A(n8302), .B(n8254), .Z(n8209) );
  HS65_LL_IVX9 U16307 ( .A(n2883), .Z(n656) );
  HS65_LL_NAND2X7 U16308 ( .A(n5472), .B(n5013), .Z(n4487) );
  HS65_LL_NAND2X7 U16309 ( .A(n7064), .B(n6606), .Z(n6080) );
  HS65_LL_NAND2X7 U16310 ( .A(n7768), .B(n7941), .Z(n8507) );
  HS65_LL_IVX9 U16311 ( .A(n3095), .Z(n213) );
  HS65_LL_NAND3X5 U16312 ( .A(n7619), .B(n7636), .C(n7637), .Z(n7635) );
  HS65_LL_NAND3X5 U16313 ( .A(n7656), .B(n7657), .C(n7658), .Z(n7655) );
  HS65_LL_NAND2X7 U16314 ( .A(n3615), .B(n2914), .Z(n3541) );
  HS65_LL_NAND3X5 U16315 ( .A(n4988), .B(n5554), .C(n4788), .Z(n5636) );
  HS65_LL_NAND3X5 U16316 ( .A(n6581), .B(n7146), .C(n6381), .Z(n7228) );
  HS65_LL_NAND3X5 U16317 ( .A(n4876), .B(n5532), .C(n4726), .Z(n5610) );
  HS65_LL_NAND3X5 U16318 ( .A(n6469), .B(n7124), .C(n6342), .Z(n7202) );
  HS65_LL_NAND3X5 U16319 ( .A(n6455), .B(n7171), .C(n6235), .Z(n7174) );
  HS65_LL_NAND3X5 U16320 ( .A(n4862), .B(n5579), .C(n4642), .Z(n5582) );
  HS65_LL_NAND3X5 U16321 ( .A(n3140), .B(n3293), .C(n3127), .Z(n4019) );
  HS65_LL_NAND2X7 U16322 ( .A(n556), .B(n6074), .Z(n6149) );
  HS65_LL_NAND2X7 U16323 ( .A(n34), .B(n4481), .Z(n4556) );
  HS65_LL_NOR2X6 U16324 ( .A(n7952), .B(n8039), .Z(n8521) );
  HS65_LL_NOR2X6 U16325 ( .A(n1985), .B(n1920), .Z(n1934) );
  HS65_LL_NOR2X6 U16326 ( .A(n4456), .B(n4448), .Z(n4758) );
  HS65_LL_NOR2X6 U16327 ( .A(n6441), .B(n6402), .Z(n6232) );
  HS65_LL_NOR2X6 U16328 ( .A(n4495), .B(n4509), .Z(n4785) );
  HS65_LL_NOR2X6 U16329 ( .A(n6088), .B(n6102), .Z(n6378) );
  HS65_LL_NOR2X6 U16330 ( .A(n6049), .B(n6041), .Z(n6339) );
  HS65_LL_NOR2X6 U16331 ( .A(n4848), .B(n4809), .Z(n4639) );
  HS65_LL_NOR2X6 U16332 ( .A(n7847), .B(n7981), .Z(n8224) );
  HS65_LL_NOR2X6 U16333 ( .A(n4549), .B(n4667), .Z(n5022) );
  HS65_LL_NOR2X6 U16334 ( .A(n6142), .B(n6260), .Z(n6615) );
  HS65_LL_IVX9 U16335 ( .A(n7064), .Z(n537) );
  HS65_LL_IVX9 U16336 ( .A(n5472), .Z(n15) );
  HS65_LL_IVX9 U16337 ( .A(n3269), .Z(n168) );
  HS65_LL_NOR2X6 U16338 ( .A(n7947), .B(n8049), .Z(n8051) );
  HS65_LL_NOR2X6 U16339 ( .A(n2361), .B(n2296), .Z(n2310) );
  HS65_LL_NOR2X6 U16340 ( .A(n3692), .B(n3342), .Z(n3705) );
  HS65_LL_IVX9 U16341 ( .A(n3157), .Z(n654) );
  HS65_LL_NOR2X6 U16342 ( .A(n2915), .B(n3047), .Z(n3644) );
  HS65_LL_NOR4ABX2 U16343 ( .A(n8849), .B(n8850), .C(n7774), .D(n8622), .Z(
        n8848) );
  HS65_LL_OA212X4 U16344 ( .A(n7768), .B(n8363), .C(n7943), .D(n8049), .E(
        n8869), .Z(n8850) );
  HS65_LL_NOR2X6 U16345 ( .A(n8150), .B(n8146), .Z(n7812) );
  HS65_LL_NOR2X6 U16346 ( .A(n8173), .B(n8169), .Z(n7910) );
  HS65_LL_IVX9 U16347 ( .A(n7920), .Z(n126) );
  HS65_LL_IVX9 U16348 ( .A(n7822), .Z(n606) );
  HS65_LL_NOR2X6 U16349 ( .A(n3807), .B(n3396), .Z(n3820) );
  HS65_LL_NOR2X6 U16350 ( .A(n1609), .B(n1544), .Z(n1558) );
  HS65_LL_NAND2X7 U16351 ( .A(n3342), .B(n2889), .Z(n3703) );
  HS65_LL_NAND2X7 U16352 ( .A(n3114), .B(n3116), .Z(n3461) );
  HS65_LL_NAND2X7 U16353 ( .A(n3396), .B(n2837), .Z(n3818) );
  HS65_LL_IVX9 U16354 ( .A(n7623), .Z(n617) );
  HS65_LL_IVX9 U16355 ( .A(n7663), .Z(n137) );
  HS65_LL_NAND2X7 U16356 ( .A(n6859), .B(n6515), .Z(n6832) );
  HS65_LL_NAND2X7 U16357 ( .A(n5267), .B(n4922), .Z(n5240) );
  HS65_LL_NAND2X7 U16358 ( .A(n5382), .B(n4975), .Z(n5355) );
  HS65_LL_NAND2X7 U16359 ( .A(n5150), .B(n4847), .Z(n5122) );
  HS65_LL_NAND2X7 U16360 ( .A(n6974), .B(n6568), .Z(n6947) );
  HS65_LL_NAND2X7 U16361 ( .A(n6742), .B(n6440), .Z(n6714) );
  HS65_LL_NAND4ABX3 U16362 ( .A(n6533), .B(n6534), .C(n6535), .D(n6536), .Z(
        n6192) );
  HS65_LL_OAI212X5 U16363 ( .A(n6544), .B(n6101), .C(n6094), .D(n6382), .E(
        n6545), .Z(n6533) );
  HS65_LL_NOR3AX2 U16364 ( .A(n6537), .B(n6538), .C(n6539), .Z(n6536) );
  HS65_LL_NAND3AX6 U16365 ( .A(n6540), .B(n6541), .C(n6542), .Z(n6534) );
  HS65_LL_NAND4ABX3 U16366 ( .A(n6480), .B(n6481), .C(n6482), .D(n6483), .Z(
        n6175) );
  HS65_LL_OAI212X5 U16367 ( .A(n6491), .B(n6040), .C(n6055), .D(n6343), .E(
        n6492), .Z(n6480) );
  HS65_LL_NOR3AX2 U16368 ( .A(n6484), .B(n6485), .C(n6486), .Z(n6483) );
  HS65_LL_NAND3AX6 U16369 ( .A(n6487), .B(n6488), .C(n6489), .Z(n6481) );
  HS65_LL_NAND4ABX3 U16370 ( .A(n4887), .B(n4888), .C(n4889), .D(n4890), .Z(
        n4582) );
  HS65_LL_OAI212X5 U16371 ( .A(n4898), .B(n4447), .C(n4462), .D(n4727), .E(
        n4899), .Z(n4887) );
  HS65_LL_NOR3AX2 U16372 ( .A(n4891), .B(n4892), .C(n4893), .Z(n4890) );
  HS65_LL_NAND3AX6 U16373 ( .A(n4894), .B(n4895), .C(n4896), .Z(n4888) );
  HS65_LL_NAND4ABX3 U16374 ( .A(n4940), .B(n4941), .C(n4942), .D(n4943), .Z(
        n4599) );
  HS65_LL_OAI212X5 U16375 ( .A(n4951), .B(n4508), .C(n4501), .D(n4789), .E(
        n4952), .Z(n4940) );
  HS65_LL_NOR3AX2 U16376 ( .A(n4944), .B(n4945), .C(n4946), .Z(n4943) );
  HS65_LL_NAND3AX6 U16377 ( .A(n4947), .B(n4948), .C(n4949), .Z(n4941) );
  HS65_LL_NAND4ABX3 U16378 ( .A(n6405), .B(n6406), .C(n6407), .D(n6408), .Z(
        n6122) );
  HS65_LL_OAI212X5 U16379 ( .A(n6416), .B(n6247), .C(n6116), .D(n6236), .E(
        n6417), .Z(n6405) );
  HS65_LL_NOR3AX2 U16380 ( .A(n6409), .B(n6410), .C(n6411), .Z(n6408) );
  HS65_LL_NAND3AX6 U16381 ( .A(n6412), .B(n6413), .C(n6414), .Z(n6406) );
  HS65_LL_NAND4ABX3 U16382 ( .A(n4812), .B(n4813), .C(n4814), .D(n4815), .Z(
        n4529) );
  HS65_LL_OAI212X5 U16383 ( .A(n4823), .B(n4654), .C(n4523), .D(n4643), .E(
        n4824), .Z(n4812) );
  HS65_LL_NOR3AX2 U16384 ( .A(n4816), .B(n4817), .C(n4818), .Z(n4815) );
  HS65_LL_NAND3AX6 U16385 ( .A(n4819), .B(n4820), .C(n4821), .Z(n4813) );
  HS65_LL_NAND2X7 U16386 ( .A(n7620), .B(n7835), .Z(n7684) );
  HS65_LL_NAND2X7 U16387 ( .A(n7660), .B(n7874), .Z(n7722) );
  HS65_LL_NOR2X6 U16388 ( .A(n5507), .B(n4667), .Z(n5104) );
  HS65_LL_NOR2X6 U16389 ( .A(n7099), .B(n6260), .Z(n6697) );
  HS65_LL_NOR2X6 U16390 ( .A(n7632), .B(n7822), .Z(n8748) );
  HS65_LL_NOR2X6 U16391 ( .A(n7652), .B(n7920), .Z(n8838) );
  HS65_LL_NOR2X6 U16392 ( .A(n7125), .B(n6475), .Z(n6918) );
  HS65_LL_NOR2X6 U16393 ( .A(n5533), .B(n4882), .Z(n5326) );
  HS65_LL_NOR2X6 U16394 ( .A(n5555), .B(n4994), .Z(n5441) );
  HS65_LL_NOR2X6 U16395 ( .A(n5571), .B(n4868), .Z(n5210) );
  HS65_LL_NOR2X6 U16396 ( .A(n7147), .B(n6587), .Z(n7033) );
  HS65_LL_NOR2X6 U16397 ( .A(n7163), .B(n6461), .Z(n6802) );
  HS65_LL_IVX9 U16398 ( .A(n2938), .Z(n226) );
  HS65_LL_NOR2X6 U16399 ( .A(n3380), .B(n3203), .Z(n3187) );
  HS65_LL_NOR2X6 U16400 ( .A(n3096), .B(n2938), .Z(n2960) );
  HS65_LL_OAI21X3 U16401 ( .A(n4670), .B(n4685), .C(n5657), .Z(n5699) );
  HS65_LL_OAI21X3 U16402 ( .A(n6263), .B(n6278), .C(n7249), .Z(n7291) );
  HS65_LL_NOR2X6 U16403 ( .A(n3224), .B(n3047), .Z(n3593) );
  HS65_LL_IVX9 U16404 ( .A(n7724), .Z(n110) );
  HS65_LL_NAND2X7 U16405 ( .A(n45), .B(n4481), .Z(n4701) );
  HS65_LL_NAND2X7 U16406 ( .A(n567), .B(n6074), .Z(n6294) );
  HS65_LL_NOR2X6 U16407 ( .A(n2957), .B(n3067), .Z(n3488) );
  HS65_LL_NAND2X7 U16408 ( .A(n120), .B(n7737), .Z(n8444) );
  HS65_LL_NOR2X6 U16409 ( .A(n5382), .B(n4773), .Z(n5384) );
  HS65_LL_NOR2X6 U16410 ( .A(n5267), .B(n4747), .Z(n5269) );
  HS65_LL_NOR2X6 U16411 ( .A(n6974), .B(n6366), .Z(n6976) );
  HS65_LL_NOR2X6 U16412 ( .A(n5150), .B(n4627), .Z(n5152) );
  HS65_LL_NOR2X6 U16413 ( .A(n6742), .B(n6220), .Z(n6744) );
  HS65_LL_NOR2X6 U16414 ( .A(n6859), .B(n6327), .Z(n6861) );
  HS65_LL_NOR2X6 U16415 ( .A(n7846), .B(n7981), .Z(n7983) );
  HS65_LL_NOR2X6 U16416 ( .A(n8123), .B(n7981), .Z(n7990) );
  HS65_LL_NAND2X7 U16417 ( .A(n7750), .B(n7859), .Z(n8204) );
  HS65_LL_NAND2X7 U16418 ( .A(n5028), .B(n4710), .Z(n5000) );
  HS65_LL_NAND2X7 U16419 ( .A(n6621), .B(n6303), .Z(n6593) );
  HS65_LL_NOR2X6 U16420 ( .A(n8150), .B(n7676), .Z(n8717) );
  HS65_LL_NAND2X7 U16421 ( .A(n524), .B(n6114), .Z(n6432) );
  HS65_LL_NAND2X7 U16422 ( .A(n700), .B(n4521), .Z(n4839) );
  HS65_LL_NOR2X6 U16423 ( .A(n4790), .B(n4976), .Z(n5454) );
  HS65_LL_NOR2X6 U16424 ( .A(n4644), .B(n4849), .Z(n5224) );
  HS65_LL_NOR2X6 U16425 ( .A(n6237), .B(n6442), .Z(n6816) );
  HS65_LL_NOR2X6 U16426 ( .A(n6383), .B(n6569), .Z(n7046) );
  HS65_LL_NOR2X6 U16427 ( .A(n4728), .B(n4923), .Z(n5339) );
  HS65_LL_NOR2X6 U16428 ( .A(n6344), .B(n6516), .Z(n6931) );
  HS65_LL_NOR2X6 U16429 ( .A(n4748), .B(n4882), .Z(n4760) );
  HS65_LL_NOR2X6 U16430 ( .A(n4774), .B(n4994), .Z(n4787) );
  HS65_LL_NOR2X6 U16431 ( .A(n4628), .B(n4868), .Z(n4641) );
  HS65_LL_NOR2X6 U16432 ( .A(n6367), .B(n6587), .Z(n6380) );
  HS65_LL_NOR2X6 U16433 ( .A(n6221), .B(n6461), .Z(n6234) );
  HS65_LL_NOR2X6 U16434 ( .A(n6328), .B(n6475), .Z(n6341) );
  HS65_LL_NAND2X7 U16435 ( .A(n602), .B(n7699), .Z(n7692) );
  HS65_LL_NAND2X7 U16436 ( .A(n122), .B(n7737), .Z(n7730) );
  HS65_LL_NOR2X6 U16437 ( .A(n2914), .B(n3034), .Z(n3556) );
  HS65_LL_IVX9 U16438 ( .A(n3286), .Z(n151) );
  HS65_LL_NAND2X7 U16439 ( .A(n551), .B(n6074), .Z(n6612) );
  HS65_LL_NAND2X7 U16440 ( .A(n29), .B(n4481), .Z(n5019) );
  HS65_LL_NAND2X7 U16441 ( .A(n615), .B(n7699), .Z(n8683) );
  HS65_LL_NAND2X7 U16442 ( .A(n135), .B(n7737), .Z(n8773) );
  HS65_LL_NAND2X7 U16443 ( .A(n2992), .B(n2830), .Z(n3819) );
  HS65_LL_NAND2X7 U16444 ( .A(n3464), .B(n2860), .Z(n3462) );
  HS65_LL_OAI21X3 U16445 ( .A(n7836), .B(n7675), .C(n8375), .Z(n8374) );
  HS65_LL_OAI21X3 U16446 ( .A(n7875), .B(n7713), .C(n8427), .Z(n8426) );
  HS65_LL_NOR2X6 U16447 ( .A(n3326), .B(n3140), .Z(n3160) );
  HS65_LL_IVX9 U16448 ( .A(n8173), .Z(n108) );
  HS65_LL_IVX9 U16449 ( .A(n8150), .Z(n588) );
  HS65_LL_AOI12X2 U16450 ( .A(n4477), .B(n4667), .C(n4668), .Z(n4663) );
  HS65_LL_AOI12X2 U16451 ( .A(n6070), .B(n6260), .C(n6261), .Z(n6256) );
  HS65_LL_OAI21X3 U16452 ( .A(n2495), .B(n2326), .C(n2555), .Z(n2554) );
  HS65_LL_OAI21X3 U16453 ( .A(n903), .B(n906), .C(n888), .Z(n2555) );
  HS65_LL_OAI21X3 U16454 ( .A(n1743), .B(n1574), .C(n1803), .Z(n1802) );
  HS65_LL_OAI21X3 U16455 ( .A(n821), .B(n824), .C(n806), .Z(n1803) );
  HS65_LL_NAND4ABX3 U16456 ( .A(n4963), .B(n4964), .C(n4965), .D(n4966), .Z(
        n4598) );
  HS65_LL_OAI222X2 U16457 ( .A(n4975), .B(n4495), .C(n4976), .D(n4774), .E(
        n4492), .F(n4509), .Z(n4964) );
  HS65_LL_NOR4ABX2 U16458 ( .A(n4967), .B(n4968), .C(n4969), .D(n4970), .Z(
        n4966) );
  HS65_LL_NAND3X5 U16459 ( .A(n4977), .B(n4978), .C(n4979), .Z(n4963) );
  HS65_LL_NAND4ABX3 U16460 ( .A(n6428), .B(n6429), .C(n6430), .D(n6431), .Z(
        n6121) );
  HS65_LL_OAI222X2 U16461 ( .A(n6440), .B(n6441), .C(n6442), .D(n6221), .E(
        n6443), .F(n6402), .Z(n6429) );
  HS65_LL_NOR4ABX2 U16462 ( .A(n6432), .B(n6433), .C(n6434), .D(n6435), .Z(
        n6431) );
  HS65_LL_NAND3X5 U16463 ( .A(n6444), .B(n6445), .C(n6446), .Z(n6428) );
  HS65_LL_NAND4ABX3 U16464 ( .A(n4835), .B(n4836), .C(n4837), .D(n4838), .Z(
        n4528) );
  HS65_LL_OAI222X2 U16465 ( .A(n4847), .B(n4848), .C(n4849), .D(n4628), .E(
        n4850), .F(n4809), .Z(n4836) );
  HS65_LL_NOR4ABX2 U16466 ( .A(n4839), .B(n4840), .C(n4841), .D(n4842), .Z(
        n4838) );
  HS65_LL_NAND3X5 U16467 ( .A(n4851), .B(n4852), .C(n4853), .Z(n4835) );
  HS65_LL_NOR2X6 U16468 ( .A(n1862), .B(n1920), .Z(n2016) );
  HS65_LL_OAI21X3 U16469 ( .A(n3807), .B(n3405), .C(n4290), .Z(n4289) );
  HS65_LL_OAI21X3 U16470 ( .A(n421), .B(n415), .C(n427), .Z(n4290) );
  HS65_LL_AOI12X2 U16471 ( .A(n4455), .B(n4460), .C(n4447), .Z(n4735) );
  HS65_LL_AOI12X2 U16472 ( .A(n4494), .B(n4499), .C(n4508), .Z(n4796) );
  HS65_LL_AOI12X2 U16473 ( .A(n6087), .B(n6092), .C(n6101), .Z(n6389) );
  HS65_LL_AOI12X2 U16474 ( .A(n6048), .B(n6053), .C(n6040), .Z(n6350) );
  HS65_LL_AOI12X2 U16475 ( .A(n6219), .B(n6118), .C(n6247), .Z(n6243) );
  HS65_LL_AOI12X2 U16476 ( .A(n4626), .B(n4525), .C(n4654), .Z(n4650) );
  HS65_LL_NAND2X7 U16477 ( .A(n2981), .B(n3326), .Z(n3714) );
  HS65_LL_NAND2X7 U16478 ( .A(n2992), .B(n3380), .Z(n3829) );
  HS65_LL_NAND2X7 U16479 ( .A(n3464), .B(n3096), .Z(n3473) );
  HS65_LL_NAND4ABX3 U16480 ( .A(n4697), .B(n4698), .C(n4699), .D(n4700), .Z(
        n4472) );
  HS65_LL_OAI222X2 U16481 ( .A(n4709), .B(n4710), .C(n4711), .D(n4551), .E(
        n4670), .F(n4712), .Z(n4698) );
  HS65_LL_NOR4ABX2 U16482 ( .A(n4705), .B(n4706), .C(n4707), .D(n4708), .Z(
        n4699) );
  HS65_LL_NOR4ABX2 U16483 ( .A(n4701), .B(n4702), .C(n4703), .D(n4704), .Z(
        n4700) );
  HS65_LL_NAND4ABX3 U16484 ( .A(n6290), .B(n6291), .C(n6292), .D(n6293), .Z(
        n6065) );
  HS65_LL_OAI222X2 U16485 ( .A(n6302), .B(n6303), .C(n6304), .D(n6144), .E(
        n6263), .F(n6305), .Z(n6291) );
  HS65_LL_NOR4ABX2 U16486 ( .A(n6298), .B(n6299), .C(n6300), .D(n6301), .Z(
        n6292) );
  HS65_LL_NOR4ABX2 U16487 ( .A(n6294), .B(n6295), .C(n6296), .D(n6297), .Z(
        n6293) );
  HS65_LL_NOR2X6 U16488 ( .A(n1575), .B(n1581), .Z(n1496) );
  HS65_LL_NOR2X6 U16489 ( .A(n2327), .B(n2333), .Z(n2248) );
  HS65_LL_IVX9 U16490 ( .A(n4847), .Z(n679) );
  HS65_LL_IVX9 U16491 ( .A(n6440), .Z(n503) );
  HS65_LL_NOR2X6 U16492 ( .A(n1951), .B(n1957), .Z(n1872) );
  HS65_LL_OAI21X3 U16493 ( .A(n4501), .B(n4509), .C(n4938), .Z(n4937) );
  HS65_LL_OAI21X3 U16494 ( .A(n4483), .B(n4670), .C(n4671), .Z(n4669) );
  HS65_LL_OAI21X3 U16495 ( .A(n6076), .B(n6263), .C(n6264), .Z(n6262) );
  HS65_LL_OAI21X3 U16496 ( .A(n6116), .B(n6402), .C(n6403), .Z(n6401) );
  HS65_LL_OAI21X3 U16497 ( .A(n4523), .B(n4809), .C(n4810), .Z(n4808) );
  HS65_LL_OAI21X3 U16498 ( .A(n3224), .B(n3225), .C(n3226), .Z(n3223) );
  HS65_LL_NOR2X6 U16499 ( .A(n2238), .B(n2296), .Z(n2392) );
  HS65_LL_OAI21X3 U16500 ( .A(n4447), .B(n4448), .C(n4449), .Z(n4446) );
  HS65_LL_OAI21X3 U16501 ( .A(n4654), .B(n4809), .C(n5687), .Z(n5761) );
  HS65_LL_OAI21X3 U16502 ( .A(n6247), .B(n6402), .C(n7279), .Z(n7353) );
  HS65_LL_OAI21X3 U16503 ( .A(n6040), .B(n6041), .C(n6042), .Z(n6039) );
  HS65_LL_NAND4ABX3 U16504 ( .A(n8404), .B(n8405), .C(n8406), .D(n8407), .Z(
        n7999) );
  HS65_LL_OAI222X2 U16505 ( .A(n7822), .B(n7620), .C(n7835), .D(n7676), .E(
        n7807), .F(n8132), .Z(n8405) );
  HS65_LL_NOR3AX2 U16506 ( .A(n8408), .B(n7792), .C(n8409), .Z(n8407) );
  HS65_LL_NOR3AX2 U16507 ( .A(n8410), .B(n8411), .C(n8412), .Z(n8406) );
  HS65_LL_NAND4ABX3 U16508 ( .A(n8456), .B(n8457), .C(n8458), .D(n8459), .Z(
        n8012) );
  HS65_LL_OAI222X2 U16509 ( .A(n7920), .B(n7660), .C(n7874), .D(n7714), .E(
        n7905), .F(n8183), .Z(n8457) );
  HS65_LL_NOR3AX2 U16510 ( .A(n8460), .B(n7891), .C(n8461), .Z(n8459) );
  HS65_LL_NOR3AX2 U16511 ( .A(n8462), .B(n8463), .C(n8464), .Z(n8458) );
  HS65_LL_NOR2X6 U16512 ( .A(n1486), .B(n1544), .Z(n1640) );
  HS65_LL_AOI12X2 U16513 ( .A(n7951), .B(n8369), .C(n7949), .Z(n8365) );
  HS65_LL_AOI12X2 U16514 ( .A(n7850), .B(n8123), .C(n7848), .Z(n8119) );
  HS65_LL_NAND2X7 U16515 ( .A(n3588), .B(n2918), .Z(n3586) );
  HS65_LL_AOI12X2 U16516 ( .A(n3032), .B(n3053), .C(n3054), .Z(n3050) );
  HS65_LL_NAND4ABX3 U16517 ( .A(n3478), .B(n3479), .C(n3480), .D(n3481), .Z(
        n2942) );
  HS65_LL_NOR3X4 U16518 ( .A(n3486), .B(n3487), .C(n3488), .Z(n3480) );
  HS65_LL_NAND4ABX3 U16519 ( .A(n3492), .B(n3493), .C(n3494), .D(n3495), .Z(
        n3478) );
  HS65_LL_OAI212X5 U16520 ( .A(n3489), .B(n3115), .C(n2857), .D(n2860), .E(
        n3490), .Z(n3479) );
  HS65_LL_NAND4ABX3 U16521 ( .A(n6728), .B(n6729), .C(n6730), .D(n6731), .Z(
        n6212) );
  HS65_LL_NOR3AX2 U16522 ( .A(n6736), .B(n6737), .C(n6738), .Z(n6730) );
  HS65_LL_OAI212X5 U16523 ( .A(n6739), .B(n6740), .C(n6462), .D(n6127), .E(
        n6741), .Z(n6729) );
  HS65_LL_NOR4ABX2 U16524 ( .A(n6732), .B(n6733), .C(n6734), .D(n6735), .Z(
        n6731) );
  HS65_LL_NAND4ABX3 U16525 ( .A(n5136), .B(n5137), .C(n5138), .D(n5139), .Z(
        n4619) );
  HS65_LL_NOR3AX2 U16526 ( .A(n5144), .B(n5145), .C(n5146), .Z(n5138) );
  HS65_LL_OAI212X5 U16527 ( .A(n5147), .B(n5148), .C(n4869), .D(n4534), .E(
        n5149), .Z(n5137) );
  HS65_LL_NOR4ABX2 U16528 ( .A(n5140), .B(n5141), .C(n5142), .D(n5143), .Z(
        n5139) );
  HS65_LL_NAND4ABX3 U16529 ( .A(n5368), .B(n5369), .C(n5370), .D(n5371), .Z(
        n4766) );
  HS65_LL_NOR3AX2 U16530 ( .A(n5376), .B(n5377), .C(n5378), .Z(n5370) );
  HS65_LL_OAI212X5 U16531 ( .A(n5379), .B(n5380), .C(n4995), .D(n4493), .E(
        n5381), .Z(n5369) );
  HS65_LL_NOR4ABX2 U16532 ( .A(n5372), .B(n5373), .C(n5374), .D(n5375), .Z(
        n5371) );
  HS65_LL_NAND4ABX3 U16533 ( .A(n6960), .B(n6961), .C(n6962), .D(n6963), .Z(
        n6359) );
  HS65_LL_NOR3AX2 U16534 ( .A(n6968), .B(n6969), .C(n6970), .Z(n6962) );
  HS65_LL_OAI212X5 U16535 ( .A(n6971), .B(n6972), .C(n6588), .D(n6086), .E(
        n6973), .Z(n6961) );
  HS65_LL_NOR4ABX2 U16536 ( .A(n6964), .B(n6965), .C(n6966), .D(n6967), .Z(
        n6963) );
  HS65_LL_AOI12X2 U16537 ( .A(n2276), .B(n2333), .C(n2274), .Z(n2329) );
  HS65_LL_AOI12X2 U16538 ( .A(n1524), .B(n1581), .C(n1522), .Z(n1577) );
  HS65_LL_AOI12X2 U16539 ( .A(n1900), .B(n1957), .C(n1898), .Z(n1953) );
  HS65_LL_AOI12X2 U16540 ( .A(n1148), .B(n1205), .C(n1146), .Z(n1201) );
  HS65_LL_NOR2X6 U16541 ( .A(n3061), .B(n3067), .Z(n3446) );
  HS65_LL_IVX9 U16542 ( .A(n3053), .Z(n142) );
  HS65_LL_NOR2X6 U16543 ( .A(n3406), .B(n3412), .Z(n2840) );
  HS65_LL_OAI21X3 U16544 ( .A(n3692), .B(n3292), .C(n4231), .Z(n4230) );
  HS65_LL_OAI21X3 U16545 ( .A(n639), .B(n633), .C(n658), .Z(n4231) );
  HS65_LL_AOI12X2 U16546 ( .A(n2917), .B(n3286), .C(n2915), .Z(n3282) );
  HS65_LL_NAND2X7 U16547 ( .A(n3588), .B(n3252), .Z(n3598) );
  HS65_LL_NOR2X6 U16548 ( .A(n7847), .B(n8649), .Z(n7968) );
  HS65_LL_NAND2X7 U16549 ( .A(n1519), .B(n1486), .Z(n1662) );
  HS65_LL_NAND2X7 U16550 ( .A(n2271), .B(n2238), .Z(n2414) );
  HS65_LL_IVX9 U16551 ( .A(n3252), .Z(n154) );
  HS65_LL_NOR2X6 U16552 ( .A(n3984), .B(n2914), .Z(n3049) );
  HS65_LL_NOR2X6 U16553 ( .A(n4571), .B(n5501), .Z(n5029) );
  HS65_LL_NOR2X6 U16554 ( .A(n6164), .B(n7093), .Z(n6622) );
  HS65_LL_NAND2X7 U16555 ( .A(n7941), .B(n8510), .Z(n7946) );
  HS65_LL_NAND2X7 U16556 ( .A(n8510), .B(n8057), .Z(n8538) );
  HS65_LL_AOI12X2 U16557 ( .A(n7686), .B(n8150), .C(n8421), .Z(n8417) );
  HS65_LL_AOI12X2 U16558 ( .A(n7724), .B(n8173), .C(n8473), .Z(n8469) );
  HS65_LL_NOR2X6 U16559 ( .A(n6742), .B(n6221), .Z(n6233) );
  HS65_LL_NOR2X6 U16560 ( .A(n5150), .B(n4628), .Z(n4640) );
  HS65_LL_NAND2X7 U16561 ( .A(n7821), .B(n7806), .Z(n8747) );
  HS65_LL_NAND2X7 U16562 ( .A(n7919), .B(n7869), .Z(n8837) );
  HS65_LL_NAND2X7 U16563 ( .A(n4593), .B(n4454), .Z(n5316) );
  HS65_LL_NAND2X7 U16564 ( .A(n4610), .B(n4493), .Z(n5431) );
  HS65_LL_NAND2X7 U16565 ( .A(n6186), .B(n6047), .Z(n6908) );
  HS65_LL_NAND2X7 U16566 ( .A(n5135), .B(n4534), .Z(n5200) );
  HS65_LL_NAND2X7 U16567 ( .A(n6203), .B(n6086), .Z(n7023) );
  HS65_LL_NAND2X7 U16568 ( .A(n6727), .B(n6127), .Z(n6792) );
  HS65_LL_NAND2X7 U16569 ( .A(n8207), .B(n7851), .Z(n8205) );
  HS65_LL_NOR2X6 U16570 ( .A(n6278), .B(n6621), .Z(n6642) );
  HS65_LL_NOR2X6 U16571 ( .A(n4685), .B(n5028), .Z(n5049) );
  HS65_LL_NAND2X7 U16572 ( .A(n2271), .B(n2361), .Z(n2429) );
  HS65_LL_NAND2X7 U16573 ( .A(n1519), .B(n1609), .Z(n1677) );
  HS65_LL_NAND2X7 U16574 ( .A(n6114), .B(n525), .Z(n6227) );
  HS65_LL_NAND2X7 U16575 ( .A(n4606), .B(n467), .Z(n4780) );
  HS65_LL_NAND2X7 U16576 ( .A(n6199), .B(n292), .Z(n6373) );
  HS65_LL_NAND2X7 U16577 ( .A(n4521), .B(n701), .Z(n4634) );
  HS65_LL_AOI12X2 U16578 ( .A(n7767), .B(n8556), .C(n8058), .Z(n8870) );
  HS65_LL_NAND2X7 U16579 ( .A(n564), .B(n6074), .Z(n6676) );
  HS65_LL_NAND2X7 U16580 ( .A(n42), .B(n4481), .Z(n5083) );
  HS65_LL_AOI12X2 U16581 ( .A(n4670), .B(n5028), .C(n5026), .Z(n5479) );
  HS65_LL_AOI12X2 U16582 ( .A(n6263), .B(n6621), .C(n6619), .Z(n7071) );
  HS65_LL_IVX9 U16583 ( .A(n3615), .Z(n158) );
  HS65_LL_NOR2X6 U16584 ( .A(n7656), .B(n8776), .Z(n8779) );
  HS65_LL_NOR2X6 U16585 ( .A(n7619), .B(n8686), .Z(n8689) );
  HS65_LL_NOR2X6 U16586 ( .A(n3225), .B(n3034), .Z(n3259) );
  HS65_LL_NAND2X7 U16587 ( .A(n7821), .B(n8155), .Z(n8674) );
  HS65_LL_NAND2X7 U16588 ( .A(n7919), .B(n8178), .Z(n8764) );
  HS65_LL_NAND2X7 U16589 ( .A(n6727), .B(n6442), .Z(n6723) );
  HS65_LL_NAND2X7 U16590 ( .A(n5135), .B(n4849), .Z(n5131) );
  HS65_LL_NAND2X7 U16591 ( .A(n6186), .B(n6516), .Z(n6841) );
  HS65_LL_NAND2X7 U16592 ( .A(n4593), .B(n4923), .Z(n5249) );
  HS65_LL_NAND2X7 U16593 ( .A(n4610), .B(n4976), .Z(n5364) );
  HS65_LL_NAND2X7 U16594 ( .A(n6203), .B(n6569), .Z(n6956) );
  HS65_LL_NOR2X6 U16595 ( .A(n4667), .B(n5026), .Z(n5108) );
  HS65_LL_NOR2X6 U16596 ( .A(n6260), .B(n6619), .Z(n6701) );
  HS65_LL_NOR2X6 U16597 ( .A(n8369), .B(n8363), .Z(n8523) );
  HS65_LL_NOR2X6 U16598 ( .A(n8123), .B(n8117), .Z(n8298) );
  HS65_LL_NAND2X7 U16599 ( .A(n7859), .B(n8207), .Z(n7864) );
  HS65_LL_NOR2X6 U16600 ( .A(n3157), .B(n3342), .Z(n3333) );
  HS65_LL_NAND2X7 U16601 ( .A(n697), .B(n4521), .Z(n5205) );
  HS65_LL_NAND2X7 U16602 ( .A(n521), .B(n6114), .Z(n6797) );
  HS65_LL_NAND2X7 U16603 ( .A(n569), .B(n6074), .Z(n6630) );
  HS65_LL_NAND2X7 U16604 ( .A(n47), .B(n4481), .Z(n5037) );
  HS65_LL_NAND2X7 U16605 ( .A(n8661), .B(n7848), .Z(n8492) );
  HS65_LL_AOI12X2 U16606 ( .A(n3225), .B(n3615), .C(n3269), .Z(n3913) );
  HS65_LL_NOR2X6 U16607 ( .A(n8145), .B(n7620), .Z(n7788) );
  HS65_LL_NOR2X6 U16608 ( .A(n8168), .B(n7660), .Z(n7887) );
  HS65_LL_AOI12X2 U16609 ( .A(n7675), .B(n8686), .C(n7822), .Z(n9050) );
  HS65_LL_AOI12X2 U16610 ( .A(n7713), .B(n8776), .C(n7920), .Z(n9108) );
  HS65_LL_IVX9 U16611 ( .A(n4849), .Z(n680) );
  HS65_LL_IVX9 U16612 ( .A(n6442), .Z(n504) );
  HS65_LL_NOR2X6 U16613 ( .A(n5533), .B(n4923), .Z(n4930) );
  HS65_LL_NOR2X6 U16614 ( .A(n5555), .B(n4976), .Z(n4983) );
  HS65_LL_NOR2X6 U16615 ( .A(n7125), .B(n6516), .Z(n6523) );
  HS65_LL_NOR2X6 U16616 ( .A(n7147), .B(n6569), .Z(n6576) );
  HS65_LL_NOR2X6 U16617 ( .A(n7163), .B(n6442), .Z(n6450) );
  HS65_LL_NOR2X6 U16618 ( .A(n5571), .B(n4849), .Z(n4857) );
  HS65_LL_NOR2X6 U16619 ( .A(n6070), .B(n6144), .Z(n6662) );
  HS65_LL_NOR2X6 U16620 ( .A(n4477), .B(n4551), .Z(n5069) );
  HS65_LL_NAND2X7 U16621 ( .A(n7699), .B(n603), .Z(n7693) );
  HS65_LL_NAND2X7 U16622 ( .A(n7737), .B(n123), .Z(n7731) );
  HS65_LL_NOR2X6 U16623 ( .A(n7980), .B(n7992), .Z(n8225) );
  HS65_LL_IVX9 U16624 ( .A(n4551), .Z(n46) );
  HS65_LL_IVX9 U16625 ( .A(n6144), .Z(n568) );
  HS65_LL_NAND2X7 U16626 ( .A(n4481), .B(n40), .Z(n4714) );
  HS65_LL_NAND2X7 U16627 ( .A(n6074), .B(n562), .Z(n6307) );
  HS65_LL_NAND3X5 U16628 ( .A(n1920), .B(n1951), .C(n1907), .Z(n2171) );
  HS65_LL_IVX9 U16629 ( .A(n3034), .Z(n179) );
  HS65_LL_NAND2X7 U16630 ( .A(n8871), .B(n7949), .Z(n8619) );
  HS65_LL_NAND3X5 U16631 ( .A(n2296), .B(n2327), .C(n2283), .Z(n2547) );
  HS65_LL_NAND2X7 U16632 ( .A(n4606), .B(n482), .Z(n4978) );
  HS65_LL_NAND2X7 U16633 ( .A(n6199), .B(n307), .Z(n6571) );
  HS65_LL_NAND2X7 U16634 ( .A(n6114), .B(n519), .Z(n6445) );
  HS65_LL_NAND2X7 U16635 ( .A(n4521), .B(n695), .Z(n4852) );
  HS65_LL_NOR2X6 U16636 ( .A(n8179), .B(n7663), .Z(n8826) );
  HS65_LL_NOR2X6 U16637 ( .A(n8128), .B(n7623), .Z(n8736) );
  HS65_LL_NOR2X6 U16638 ( .A(n6126), .B(n6221), .Z(n6783) );
  HS65_LL_NOR2X6 U16639 ( .A(n4533), .B(n4628), .Z(n5191) );
  HS65_LL_NOR2X6 U16640 ( .A(n6179), .B(n6328), .Z(n6899) );
  HS65_LL_NOR2X6 U16641 ( .A(n4586), .B(n4748), .Z(n5307) );
  HS65_LL_NOR2X6 U16642 ( .A(n4603), .B(n4774), .Z(n5422) );
  HS65_LL_NOR2X6 U16643 ( .A(n6196), .B(n6367), .Z(n7014) );
  HS65_LL_NOR2X6 U16644 ( .A(n4847), .B(n4627), .Z(n5214) );
  HS65_LL_NOR2X6 U16645 ( .A(n6440), .B(n6220), .Z(n6806) );
  HS65_LL_NAND3X5 U16646 ( .A(n1544), .B(n1575), .C(n1531), .Z(n1795) );
  HS65_LL_NAND2X7 U16647 ( .A(n510), .B(n6114), .Z(n6733) );
  HS65_LL_NAND2X7 U16648 ( .A(n686), .B(n4521), .Z(n5141) );
  HS65_LL_OAI21X3 U16649 ( .A(n2119), .B(n1950), .C(n2179), .Z(n2178) );
  HS65_LL_OAI21X3 U16650 ( .A(n780), .B(n783), .C(n765), .Z(n2179) );
  HS65_LL_IVX9 U16651 ( .A(n4748), .Z(n250) );
  HS65_LL_IVX9 U16652 ( .A(n4774), .Z(n467) );
  HS65_LL_IVX9 U16653 ( .A(n4628), .Z(n701) );
  HS65_LL_IVX9 U16654 ( .A(n6367), .Z(n292) );
  HS65_LL_IVX9 U16655 ( .A(n6221), .Z(n525) );
  HS65_LL_CBI4I1X5 U16656 ( .A(n1520), .B(n1521), .C(n1522), .D(n1523), .Z(
        n1510) );
  HS65_LL_OAI21X3 U16657 ( .A(n799), .B(n814), .C(n827), .Z(n1523) );
  HS65_LL_NAND2X7 U16658 ( .A(n526), .B(n6114), .Z(n6751) );
  HS65_LL_NAND2X7 U16659 ( .A(n702), .B(n4521), .Z(n5159) );
  HS65_LL_NAND2X7 U16660 ( .A(n469), .B(n4606), .Z(n5391) );
  HS65_LL_NAND2X7 U16661 ( .A(n294), .B(n6199), .Z(n6983) );
  HS65_LL_NAND2X7 U16662 ( .A(n5013), .B(n4478), .Z(n5078) );
  HS65_LL_NAND2X7 U16663 ( .A(n6606), .B(n6071), .Z(n6671) );
  HS65_LL_NAND3X5 U16664 ( .A(n2938), .B(n3061), .C(n2925), .Z(n3929) );
  HS65_LL_NAND3X5 U16665 ( .A(n3203), .B(n3406), .C(n3191), .Z(n4042) );
  HS65_LL_AOI12X2 U16666 ( .A(n1544), .B(n1545), .C(n1505), .Z(n1540) );
  HS65_LL_AOI12X2 U16667 ( .A(n2296), .B(n2297), .C(n2257), .Z(n2292) );
  HS65_LL_AOI12X2 U16668 ( .A(n1920), .B(n1921), .C(n1881), .Z(n1916) );
  HS65_LL_AOI12X2 U16669 ( .A(n1168), .B(n1169), .C(n1129), .Z(n1164) );
  HS65_LL_NAND3X5 U16670 ( .A(n7942), .B(n8363), .C(n8027), .Z(n8933) );
  HS65_LL_NAND3X5 U16671 ( .A(n7860), .B(n8117), .C(n7959), .Z(n8993) );
  HS65_LL_NAND4ABX3 U16672 ( .A(n8388), .B(n8389), .C(n8390), .D(n8391), .Z(
        n7998) );
  HS65_LL_OAI222X2 U16673 ( .A(n8397), .B(n7831), .C(n8146), .D(n8155), .E(
        n7676), .F(n7675), .Z(n8389) );
  HS65_LL_NOR4ABX2 U16674 ( .A(n8394), .B(n8395), .C(n8396), .D(n7825), .Z(
        n8390) );
  HS65_LL_NAND3AX6 U16675 ( .A(n7813), .B(n8398), .C(n8399), .Z(n8388) );
  HS65_LL_NAND4ABX3 U16676 ( .A(n8440), .B(n8441), .C(n8442), .D(n8443), .Z(
        n8011) );
  HS65_LL_OAI222X2 U16677 ( .A(n8449), .B(n7870), .C(n8169), .D(n8178), .E(
        n7714), .F(n7713), .Z(n8441) );
  HS65_LL_NOR4ABX2 U16678 ( .A(n8446), .B(n8447), .C(n8448), .D(n7923), .Z(
        n8442) );
  HS65_LL_NAND3AX6 U16679 ( .A(n7911), .B(n8450), .C(n8451), .Z(n8440) );
  HS65_LL_NAND2X7 U16680 ( .A(n131), .B(n7737), .Z(n8447) );
  HS65_LL_NAND2X7 U16681 ( .A(n611), .B(n7699), .Z(n8395) );
  HS65_LL_IVX9 U16682 ( .A(n4711), .Z(n25) );
  HS65_LL_IVX9 U16683 ( .A(n6304), .Z(n547) );
  HS65_LL_NAND2X7 U16684 ( .A(n6606), .B(n6304), .Z(n6602) );
  HS65_LL_NAND2X7 U16685 ( .A(n5013), .B(n4711), .Z(n5009) );
  HS65_LL_AOI12X2 U16686 ( .A(n3203), .B(n3204), .C(n2845), .Z(n3199) );
  HS65_LL_AOI12X2 U16687 ( .A(n3140), .B(n3141), .C(n2875), .Z(n3136) );
  HS65_LL_NOR2X6 U16688 ( .A(n2957), .B(n2859), .Z(n3434) );
  HS65_LL_NOR2X6 U16689 ( .A(n3183), .B(n2997), .Z(n3792) );
  HS65_LL_NOR2X6 U16690 ( .A(n3157), .B(n2972), .Z(n3677) );
  HS65_LL_AOI12X2 U16691 ( .A(n7942), .B(n8039), .C(n7767), .Z(n8035) );
  HS65_LL_NOR4ABX2 U16692 ( .A(n8483), .B(n8484), .C(n7756), .D(n8485), .Z(
        n8478) );
  HS65_LL_OA212X4 U16693 ( .A(n7750), .B(n8117), .C(n7861), .D(n7981), .E(
        n8491), .Z(n8484) );
  HS65_LL_AOI12X2 U16694 ( .A(n2938), .B(n2939), .C(n2940), .Z(n2934) );
  HS65_LL_AOI12X2 U16695 ( .A(n7860), .B(n7971), .C(n7749), .Z(n7967) );
  HS65_LL_NAND4ABX3 U16696 ( .A(n3239), .B(n3240), .C(n3241), .D(n3242), .Z(
        n2910) );
  HS65_LL_OAI222X2 U16697 ( .A(n3251), .B(n2914), .C(n3034), .D(n3252), .E(
        n3253), .F(n3225), .Z(n3240) );
  HS65_LL_NAND3AX6 U16698 ( .A(n3254), .B(n3255), .C(n3256), .Z(n3239) );
  HS65_LL_NOR4ABX2 U16699 ( .A(n3243), .B(n3244), .C(n3245), .D(n3246), .Z(
        n3242) );
  HS65_LL_NOR2X6 U16700 ( .A(n3286), .B(n3034), .Z(n3037) );
  HS65_LL_NAND4ABX3 U16701 ( .A(n3083), .B(n3084), .C(n3085), .D(n3086), .Z(
        n2867) );
  HS65_LL_OAI222X2 U16702 ( .A(n3095), .B(n2856), .C(n2958), .D(n3096), .E(
        n2940), .F(n3097), .Z(n3084) );
  HS65_LL_NOR4ABX2 U16703 ( .A(n3091), .B(n3092), .C(n3093), .D(n3094), .Z(
        n3085) );
  HS65_LL_NOR4ABX2 U16704 ( .A(n3087), .B(n3088), .C(n3089), .D(n3090), .Z(
        n3086) );
  HS65_LL_NAND4ABX3 U16705 ( .A(n3368), .B(n3369), .C(n3370), .D(n3371), .Z(
        n2990) );
  HS65_LL_OAI222X2 U16706 ( .A(n2831), .B(n2994), .C(n3185), .D(n3380), .E(
        n2845), .F(n2829), .Z(n3369) );
  HS65_LL_NOR4ABX2 U16707 ( .A(n3376), .B(n3377), .C(n3378), .D(n3379), .Z(
        n3370) );
  HS65_LL_NOR4ABX2 U16708 ( .A(n3372), .B(n3373), .C(n3374), .D(n3375), .Z(
        n3371) );
  HS65_LL_IVX9 U16709 ( .A(n4534), .Z(n678) );
  HS65_LL_NAND2X7 U16710 ( .A(n6074), .B(n568), .Z(n6150) );
  HS65_LL_NAND2X7 U16711 ( .A(n4481), .B(n46), .Z(n4557) );
  HS65_LL_NAND2X7 U16712 ( .A(n4606), .B(n474), .Z(n4971) );
  HS65_LL_NAND2X7 U16713 ( .A(n6199), .B(n299), .Z(n6564) );
  HS65_LL_NAND2X7 U16714 ( .A(n4521), .B(n688), .Z(n4843) );
  HS65_LL_NAND2X7 U16715 ( .A(n6114), .B(n512), .Z(n6436) );
  HS65_LL_IVX9 U16716 ( .A(n5028), .Z(n20) );
  HS65_LL_IVX9 U16717 ( .A(n6621), .Z(n542) );
  HS65_LL_AOI12X2 U16718 ( .A(n8058), .B(n8630), .C(n7941), .Z(n8868) );
  HS65_LL_AOI12X2 U16719 ( .A(n5026), .B(n5514), .C(n5472), .Z(n5650) );
  HS65_LL_AOI12X2 U16720 ( .A(n6619), .B(n7106), .C(n7064), .Z(n7242) );
  HS65_LL_NOR2X6 U16721 ( .A(n7713), .B(n8168), .Z(n7911) );
  HS65_LL_NOR2X6 U16722 ( .A(n7675), .B(n8145), .Z(n7813) );
  HS65_LL_IVX9 U16723 ( .A(n4667), .Z(n22) );
  HS65_LL_IVX9 U16724 ( .A(n6260), .Z(n544) );
  HS65_LL_AOI12X2 U16725 ( .A(n348), .B(n7946), .C(n8616), .Z(n8615) );
  HS65_LL_AOI12X2 U16726 ( .A(n8540), .B(n7941), .C(n8313), .Z(n8616) );
  HS65_LL_AOI12X2 U16727 ( .A(n387), .B(n7864), .C(n8658), .Z(n8657) );
  HS65_LL_AOI12X2 U16728 ( .A(n8238), .B(n7859), .C(n8067), .Z(n8658) );
  HS65_LL_IVX9 U16729 ( .A(n5382), .Z(n455) );
  HS65_LL_IVX9 U16730 ( .A(n5150), .Z(n675) );
  HS65_LL_IVX9 U16731 ( .A(n6742), .Z(n499) );
  HS65_LL_AOI12X2 U16732 ( .A(n2859), .B(n3067), .C(n2857), .Z(n3063) );
  HS65_LL_AOI12X2 U16733 ( .A(n2972), .B(n3299), .C(n2970), .Z(n3295) );
  HS65_LL_AOI12X2 U16734 ( .A(n2997), .B(n3412), .C(n2995), .Z(n3408) );
  HS65_LL_AOI12X2 U16735 ( .A(n843), .B(n1114), .C(n1115), .Z(n1113) );
  HS65_LL_AOI12X2 U16736 ( .A(n1116), .B(n1117), .C(n1118), .Z(n1115) );
  HS65_LL_AOI12X2 U16737 ( .A(n761), .B(n1866), .C(n1867), .Z(n1865) );
  HS65_LL_AOI12X2 U16738 ( .A(n1868), .B(n1869), .C(n1870), .Z(n1867) );
  HS65_LL_AOI12X2 U16739 ( .A(n884), .B(n2242), .C(n2243), .Z(n2241) );
  HS65_LL_AOI12X2 U16740 ( .A(n2244), .B(n2245), .C(n2246), .Z(n2243) );
  HS65_LL_AOI12X2 U16741 ( .A(n802), .B(n1490), .C(n1491), .Z(n1489) );
  HS65_LL_AOI12X2 U16742 ( .A(n1492), .B(n1493), .C(n1494), .Z(n1491) );
  HS65_LL_AOI12X2 U16743 ( .A(n431), .B(n2834), .C(n2835), .Z(n2833) );
  HS65_LL_AOI12X2 U16744 ( .A(n2836), .B(n2837), .C(n2838), .Z(n2835) );
  HS65_LL_AOI12X2 U16745 ( .A(n225), .B(n2869), .C(n4223), .Z(n4222) );
  HS65_LL_AOI12X2 U16746 ( .A(n3475), .B(n3116), .C(n3069), .Z(n4223) );
  HS65_LL_AOI12X2 U16747 ( .A(n644), .B(n2886), .C(n2887), .Z(n2885) );
  HS65_LL_AOI12X2 U16748 ( .A(n2888), .B(n2889), .C(n2890), .Z(n2887) );
  HS65_LL_AOI12X2 U16749 ( .A(n178), .B(n3045), .C(n3046), .Z(n3044) );
  HS65_LL_AOI12X2 U16750 ( .A(n3047), .B(n3035), .C(n3048), .Z(n3046) );
  HS65_LL_AOI12X2 U16751 ( .A(n45), .B(n4569), .C(n4570), .Z(n4568) );
  HS65_LL_AOI12X2 U16752 ( .A(n4571), .B(n4552), .C(n4572), .Z(n4570) );
  HS65_LL_AOI12X2 U16753 ( .A(n567), .B(n6162), .C(n6163), .Z(n6161) );
  HS65_LL_AOI12X2 U16754 ( .A(n6164), .B(n6145), .C(n6165), .Z(n6163) );
  HS65_LL_AOI12X2 U16755 ( .A(n600), .B(n8130), .C(n8131), .Z(n8129) );
  HS65_LL_AOI12X2 U16756 ( .A(n8132), .B(n7624), .C(n7622), .Z(n8131) );
  HS65_LL_AOI12X2 U16757 ( .A(n120), .B(n8181), .C(n8182), .Z(n8180) );
  HS65_LL_AOI12X2 U16758 ( .A(n8183), .B(n7664), .C(n7662), .Z(n8182) );
  HS65_LL_AOI12X2 U16759 ( .A(n646), .B(n3131), .C(n3132), .Z(n3130) );
  HS65_LL_AOI12X2 U16760 ( .A(n3133), .B(n3134), .C(n3135), .Z(n3132) );
  HS65_LL_AOI12X2 U16761 ( .A(n253), .B(n4730), .C(n4731), .Z(n4729) );
  HS65_LL_AOI12X2 U16762 ( .A(n4732), .B(n4733), .C(n4734), .Z(n4731) );
  HS65_LL_AOI12X2 U16763 ( .A(n470), .B(n4792), .C(n4793), .Z(n4791) );
  HS65_LL_AOI12X2 U16764 ( .A(n4794), .B(n4775), .C(n4795), .Z(n4793) );
  HS65_LL_AOI12X2 U16765 ( .A(n295), .B(n6385), .C(n6386), .Z(n6384) );
  HS65_LL_AOI12X2 U16766 ( .A(n6387), .B(n6368), .C(n6388), .Z(n6386) );
  HS65_LL_AOI12X2 U16767 ( .A(n88), .B(n6346), .C(n6347), .Z(n6345) );
  HS65_LL_AOI12X2 U16768 ( .A(n6348), .B(n6329), .C(n6349), .Z(n6347) );
  HS65_LL_AOI12X2 U16769 ( .A(n524), .B(n6239), .C(n6240), .Z(n6238) );
  HS65_LL_AOI12X2 U16770 ( .A(n6241), .B(n6222), .C(n6242), .Z(n6240) );
  HS65_LL_AOI12X2 U16771 ( .A(n700), .B(n4646), .C(n4647), .Z(n4645) );
  HS65_LL_AOI12X2 U16772 ( .A(n4648), .B(n4629), .C(n4649), .Z(n4647) );
  HS65_LL_AOI12X2 U16773 ( .A(n6196), .B(n6587), .C(n6588), .Z(n6583) );
  HS65_LL_AOI12X2 U16774 ( .A(n6179), .B(n6475), .C(n6476), .Z(n6471) );
  HS65_LL_AOI12X2 U16775 ( .A(n4586), .B(n4882), .C(n4883), .Z(n4878) );
  HS65_LL_AOI12X2 U16776 ( .A(n4603), .B(n4994), .C(n4995), .Z(n4990) );
  HS65_LL_AOI12X2 U16777 ( .A(n6126), .B(n6461), .C(n6462), .Z(n6457) );
  HS65_LL_AOI12X2 U16778 ( .A(n4533), .B(n4868), .C(n4869), .Z(n4864) );
  HS65_LL_IVX9 U16779 ( .A(n6461), .Z(n501) );
  HS65_LL_IVX9 U16780 ( .A(n4868), .Z(n677) );
  HS65_LL_AOI12X2 U16781 ( .A(n467), .B(n4497), .C(n4498), .Z(n4496) );
  HS65_LL_AOI12X2 U16782 ( .A(n4499), .B(n4500), .C(n4501), .Z(n4498) );
  HS65_LL_AOI12X2 U16783 ( .A(n250), .B(n4458), .C(n4459), .Z(n4457) );
  HS65_LL_AOI12X2 U16784 ( .A(n4460), .B(n4461), .C(n4462), .Z(n4459) );
  HS65_LL_AOI12X2 U16785 ( .A(n292), .B(n6090), .C(n6091), .Z(n6089) );
  HS65_LL_AOI12X2 U16786 ( .A(n6092), .B(n6093), .C(n6094), .Z(n6091) );
  HS65_LL_AOI12X2 U16787 ( .A(n701), .B(n4527), .C(n5816), .Z(n5815) );
  HS65_LL_AOI12X2 U16788 ( .A(n4525), .B(n5496), .C(n4523), .Z(n5816) );
  HS65_LL_AOI12X2 U16789 ( .A(n525), .B(n6120), .C(n7408), .Z(n7407) );
  HS65_LL_AOI12X2 U16790 ( .A(n6118), .B(n7088), .C(n6116), .Z(n7408) );
  HS65_LL_AOI12X2 U16791 ( .A(n91), .B(n6051), .C(n6052), .Z(n6050) );
  HS65_LL_AOI12X2 U16792 ( .A(n6053), .B(n6054), .C(n6055), .Z(n6052) );
  HS65_LL_AOI12X2 U16793 ( .A(n384), .B(n7963), .C(n7964), .Z(n7962) );
  HS65_LL_AOI12X2 U16794 ( .A(n7965), .B(n7966), .C(n7858), .Z(n7964) );
  HS65_LL_AOI12X2 U16795 ( .A(n345), .B(n8031), .C(n8032), .Z(n8030) );
  HS65_LL_AOI12X2 U16796 ( .A(n8033), .B(n8034), .C(n7940), .Z(n8032) );
  HS65_LL_AOI12X2 U16797 ( .A(n123), .B(n7872), .C(n7873), .Z(n7871) );
  HS65_LL_AOI12X2 U16798 ( .A(n7652), .B(n7874), .C(n7875), .Z(n7873) );
  HS65_LL_AOI12X2 U16799 ( .A(n603), .B(n7833), .C(n7834), .Z(n7832) );
  HS65_LL_AOI12X2 U16800 ( .A(n7632), .B(n7835), .C(n7836), .Z(n7834) );
  HS65_LL_NAND2X7 U16801 ( .A(n8510), .B(n7952), .Z(n8508) );
  HS65_LL_AOI12X2 U16802 ( .A(n757), .B(n1911), .C(n1912), .Z(n1910) );
  HS65_LL_AOI12X2 U16803 ( .A(n1913), .B(n1914), .C(n1915), .Z(n1912) );
  HS65_LL_AOI12X2 U16804 ( .A(n798), .B(n1535), .C(n1536), .Z(n1534) );
  HS65_LL_AOI12X2 U16805 ( .A(n1537), .B(n1538), .C(n1539), .Z(n1536) );
  HS65_LL_AOI12X2 U16806 ( .A(n880), .B(n2287), .C(n2288), .Z(n2286) );
  HS65_LL_AOI12X2 U16807 ( .A(n2289), .B(n2290), .C(n2291), .Z(n2288) );
  HS65_LL_AOI12X2 U16808 ( .A(n433), .B(n3195), .C(n3196), .Z(n3194) );
  HS65_LL_AOI12X2 U16809 ( .A(n3197), .B(n3184), .C(n3198), .Z(n3196) );
  HS65_LL_AOI12X2 U16810 ( .A(n224), .B(n2929), .C(n2930), .Z(n2928) );
  HS65_LL_AOI12X2 U16811 ( .A(n2931), .B(n2932), .C(n2933), .Z(n2930) );
  HS65_LL_AOI12X2 U16812 ( .A(n46), .B(n4487), .C(n5754), .Z(n5753) );
  HS65_LL_AOI12X2 U16813 ( .A(n4485), .B(n5472), .C(n4483), .Z(n5754) );
  HS65_LL_AOI12X2 U16814 ( .A(n568), .B(n6080), .C(n7346), .Z(n7345) );
  HS65_LL_AOI12X2 U16815 ( .A(n6078), .B(n7064), .C(n6076), .Z(n7346) );
  HS65_LL_AOI12X2 U16816 ( .A(n179), .B(n2912), .C(n4161), .Z(n4160) );
  HS65_LL_AOI12X2 U16817 ( .A(n3053), .B(n3271), .C(n3224), .Z(n4161) );
  HS65_LL_NAND2X7 U16818 ( .A(n4481), .B(n33), .Z(n4705) );
  HS65_LL_NAND2X7 U16819 ( .A(n6074), .B(n555), .Z(n6298) );
  HS65_LL_AOI12X2 U16820 ( .A(n175), .B(n144), .C(n4079), .Z(n4078) );
  HS65_LL_AOI12X2 U16821 ( .A(n3225), .B(n3270), .C(n3253), .Z(n4079) );
  HS65_LL_IVX9 U16822 ( .A(n3279), .Z(n144) );
  HS65_LL_AOI12X2 U16823 ( .A(n264), .B(n239), .C(n5824), .Z(n5823) );
  HS65_LL_AOI12X2 U16824 ( .A(n4448), .B(n5588), .C(n4453), .Z(n5824) );
  HS65_LL_IVX9 U16825 ( .A(n4875), .Z(n239) );
  HS65_LL_AOI12X2 U16826 ( .A(n481), .B(n456), .C(n5883), .Z(n5882) );
  HS65_LL_AOI12X2 U16827 ( .A(n4509), .B(n5630), .C(n4492), .Z(n5883) );
  HS65_LL_IVX9 U16828 ( .A(n4987), .Z(n456) );
  HS65_LL_AOI12X2 U16829 ( .A(n697), .B(n667), .C(n5673), .Z(n5672) );
  HS65_LL_AOI12X2 U16830 ( .A(n4809), .B(n5581), .C(n4850), .Z(n5673) );
  HS65_LL_IVX9 U16831 ( .A(n4861), .Z(n667) );
  HS65_LL_AOI12X2 U16832 ( .A(n78), .B(n61), .C(n7416), .Z(n7415) );
  HS65_LL_AOI12X2 U16833 ( .A(n6041), .B(n7180), .C(n6046), .Z(n7416) );
  HS65_LL_IVX9 U16834 ( .A(n6468), .Z(n61) );
  HS65_LL_AOI12X2 U16835 ( .A(n306), .B(n281), .C(n7475), .Z(n7474) );
  HS65_LL_AOI12X2 U16836 ( .A(n6102), .B(n7222), .C(n6085), .Z(n7475) );
  HS65_LL_IVX9 U16837 ( .A(n6580), .Z(n281) );
  HS65_LL_AOI12X2 U16838 ( .A(n521), .B(n491), .C(n7265), .Z(n7264) );
  HS65_LL_AOI12X2 U16839 ( .A(n6402), .B(n7173), .C(n6443), .Z(n7265) );
  HS65_LL_IVX9 U16840 ( .A(n6454), .Z(n491) );
  HS65_LL_AOI12X2 U16841 ( .A(n392), .B(n364), .C(n7748), .Z(n7745) );
  HS65_LL_AOI12X2 U16842 ( .A(n7749), .B(n7750), .C(n7751), .Z(n7748) );
  HS65_LL_IVX9 U16843 ( .A(n7752), .Z(n364) );
  HS65_LL_AOI12X2 U16844 ( .A(n612), .B(n581), .C(n7674), .Z(n7671) );
  HS65_LL_AOI12X2 U16845 ( .A(n7675), .B(n7620), .C(n7676), .Z(n7674) );
  HS65_LL_IVX9 U16846 ( .A(n7677), .Z(n581) );
  HS65_LL_AOI12X2 U16847 ( .A(n132), .B(n101), .C(n7712), .Z(n7709) );
  HS65_LL_AOI12X2 U16848 ( .A(n7713), .B(n7660), .C(n7714), .Z(n7712) );
  HS65_LL_IVX9 U16849 ( .A(n7715), .Z(n101) );
  HS65_LL_NAND2X7 U16850 ( .A(n8207), .B(n7992), .Z(n8236) );
  HS65_LL_IVX9 U16851 ( .A(\u0/r0/N79 ), .Z(n706) );
  HS65_LL_AND2X4 U16852 ( .A(n7737), .B(n134), .Z(n7923) );
  HS65_LL_AND2X4 U16853 ( .A(n7699), .B(n614), .Z(n7825) );
  HS65_LL_AND2X4 U16854 ( .A(n6074), .B(n553), .Z(n6614) );
  HS65_LL_AND2X4 U16855 ( .A(n4481), .B(n31), .Z(n5021) );
  HS65_LL_BFX9 U16856 ( .A(n9143), .Z(n9148) );
  HS65_LL_MX41X7 U16857 ( .D0(n105), .S0(n122), .D1(n136), .S1(n113), .D2(n125), .S2(n7737), .D3(n108), .S3(n132), .Z(n8833) );
  HS65_LL_AND2X4 U16858 ( .A(n7737), .B(n124), .Z(n8174) );
  HS65_LL_CB4I1X9 U16859 ( .A(n3952), .B(n3141), .C(n3731), .D(n3694), .Z(
        n4018) );
  HS65_LL_CB4I1X9 U16860 ( .A(n8871), .B(n8039), .C(n8556), .D(n8529), .Z(
        n8927) );
  HS65_LL_CB4I1X9 U16861 ( .A(n8661), .B(n7971), .C(n8254), .D(n8304), .Z(
        n8976) );
  HS65_LL_AND2X4 U16862 ( .A(n7699), .B(n617), .Z(n7691) );
  HS65_LL_AND2X4 U16863 ( .A(n7737), .B(n137), .Z(n7729) );
  HS65_LL_AOI12X2 U16864 ( .A(n343), .B(n318), .C(n7766), .Z(n7763) );
  HS65_LL_AOI12X2 U16865 ( .A(n7767), .B(n7768), .C(n7769), .Z(n7766) );
  HS65_LL_IVX9 U16866 ( .A(n7770), .Z(n318) );
  HS65_LL_AOI212X4 U16867 ( .A(n14), .B(n32), .C(n42), .D(n5111), .E(n5112), 
        .Z(n5101) );
  HS65_LL_NAND2X7 U16868 ( .A(n4477), .B(n4711), .Z(n5111) );
  HS65_LL_IVX9 U16869 ( .A(n5113), .Z(n32) );
  HS65_LL_AOI212X4 U16870 ( .A(n536), .B(n554), .C(n564), .D(n6704), .E(n6705), 
        .Z(n6694) );
  HS65_LL_NAND2X7 U16871 ( .A(n6070), .B(n6304), .Z(n6704) );
  HS65_LL_IVX9 U16872 ( .A(n6706), .Z(n554) );
  HS65_LL_BFX9 U16873 ( .A(n9135), .Z(n9134) );
  HS65_LL_BFX9 U16874 ( .A(n9135), .Z(n9133) );
  HS65_LL_AND2X4 U16875 ( .A(n6114), .B(n513), .Z(n6225) );
  HS65_LL_AND2X4 U16876 ( .A(n4521), .B(n689), .Z(n4632) );
  HS65_LL_NOR2X6 U16877 ( .A(n920), .B(n919), .Z(n2596) );
  HS65_LL_NOR2X6 U16878 ( .A(n838), .B(n837), .Z(n1844) );
  HS65_LL_NOR2X6 U16879 ( .A(n797), .B(n796), .Z(n2220) );
  HS65_LL_NOR2X6 U16880 ( .A(n879), .B(n878), .Z(n1468) );
  HS65_LL_NOR2X6 U16881 ( .A(n414), .B(n423), .Z(n4330) );
  HS65_LL_NAND2X7 U16882 ( .A(n1458), .B(n1474), .Z(n1116) );
  HS65_LL_NAND2X7 U16883 ( .A(n2210), .B(n2226), .Z(n1868) );
  HS65_LL_NAND2X7 U16884 ( .A(n8929), .B(n8926), .Z(n7951) );
  HS65_LL_NAND2X7 U16885 ( .A(n8978), .B(n8979), .Z(n7850) );
  HS65_LL_NAND2X7 U16886 ( .A(n1834), .B(n1850), .Z(n1492) );
  HS65_LL_NAND2X7 U16887 ( .A(n2586), .B(n2602), .Z(n2244) );
  HS65_LL_NAND2X7 U16888 ( .A(n8917), .B(n8924), .Z(n8339) );
  HS65_LL_NAND2X7 U16889 ( .A(n4217), .B(n4201), .Z(n3475) );
  HS65_LL_NAND2X7 U16890 ( .A(n4151), .B(n4138), .Z(n3035) );
  HS65_LL_NAND2X7 U16891 ( .A(n2592), .B(n2593), .Z(n2276) );
  HS65_LL_NAND2X7 U16892 ( .A(n1840), .B(n1841), .Z(n1524) );
  HS65_LL_NAND2X7 U16893 ( .A(n2216), .B(n2217), .Z(n1900) );
  HS65_LL_NAND2X7 U16894 ( .A(n1464), .B(n1465), .Z(n1148) );
  HS65_LL_NAND2X7 U16895 ( .A(n8984), .B(n8971), .Z(n7751) );
  HS65_LL_NAND2X7 U16896 ( .A(n4140), .B(n4150), .Z(n2913) );
  HS65_LL_NAND2X7 U16897 ( .A(n4280), .B(n4277), .Z(n3133) );
  HS65_LL_NAND2X7 U16898 ( .A(n4216), .B(n4215), .Z(n3069) );
  HS65_LL_NAND2X7 U16899 ( .A(n4325), .B(n4331), .Z(n2838) );
  HS65_LL_NAND2X7 U16900 ( .A(n4157), .B(n4153), .Z(n3280) );
  HS65_LL_NAND2X7 U16901 ( .A(n8971), .B(n8992), .Z(n7993) );
  HS65_LL_NAND2X7 U16902 ( .A(n5934), .B(n5922), .Z(n5630) );
  HS65_LL_NAND2X7 U16903 ( .A(n7526), .B(n7514), .Z(n7222) );
  HS65_LL_NAND2X7 U16904 ( .A(n5875), .B(n5863), .Z(n5588) );
  HS65_LL_NAND2X7 U16905 ( .A(n7468), .B(n7457), .Z(n7180) );
  HS65_LL_NAND2X7 U16906 ( .A(n7399), .B(n7394), .Z(n7173) );
  HS65_LL_NAND2X7 U16907 ( .A(n5807), .B(n5802), .Z(n5581) );
  HS65_LL_NAND2X7 U16908 ( .A(n9043), .B(n9034), .Z(n8397) );
  HS65_LL_NAND2X7 U16909 ( .A(n9101), .B(n9092), .Z(n8449) );
  HS65_LL_NAND2X7 U16910 ( .A(n8990), .B(n8968), .Z(n7965) );
  HS65_LL_NAND2X7 U16911 ( .A(n5750), .B(n5747), .Z(n4661) );
  HS65_LL_NAND2X7 U16912 ( .A(n7342), .B(n7339), .Z(n6254) );
  HS65_LL_NAND2X7 U16913 ( .A(n8984), .B(n8991), .Z(n8082) );
  HS65_LL_NAND2X7 U16914 ( .A(n5870), .B(n5862), .Z(n5265) );
  HS65_LL_NAND2X7 U16915 ( .A(n5929), .B(n5921), .Z(n5380) );
  HS65_LL_NAND2X7 U16916 ( .A(n7453), .B(n7455), .Z(n6857) );
  HS65_LL_NAND2X7 U16917 ( .A(n7521), .B(n7513), .Z(n6972) );
  HS65_LL_NAND2X7 U16918 ( .A(n7397), .B(n7381), .Z(n6740) );
  HS65_LL_NAND2X7 U16919 ( .A(n8919), .B(n8908), .Z(n8033) );
  HS65_LL_NAND2X7 U16920 ( .A(n4265), .B(n4283), .Z(n3293) );
  HS65_LL_NAND2X7 U16921 ( .A(n9045), .B(n9027), .Z(n7636) );
  HS65_LL_NAND2X7 U16922 ( .A(n9103), .B(n9085), .Z(n7657) );
  HS65_LL_NAND2X7 U16923 ( .A(n2582), .B(n2603), .Z(n2258) );
  HS65_LL_NOR2X6 U16924 ( .A(n857), .B(n856), .Z(n1455) );
  HS65_LL_NOR2X6 U16925 ( .A(n898), .B(n897), .Z(n2583) );
  HS65_LL_NOR2X6 U16926 ( .A(n816), .B(n815), .Z(n1831) );
  HS65_LL_NAND2X7 U16927 ( .A(n4216), .B(n4219), .Z(n3450) );
  HS65_LL_NAND2X7 U16928 ( .A(n2206), .B(n2227), .Z(n1882) );
  HS65_LL_NAND2X7 U16929 ( .A(n1454), .B(n1475), .Z(n1130) );
  HS65_LL_NOR2X6 U16930 ( .A(n775), .B(n774), .Z(n2207) );
  HS65_LL_NAND2X7 U16931 ( .A(n1830), .B(n1851), .Z(n1506) );
  HS65_LL_NAND2X7 U16932 ( .A(n4211), .B(n4218), .Z(n3464) );
  HS65_LL_NAND2X7 U16933 ( .A(n4326), .B(n4342), .Z(n2992) );
  HS65_LL_NAND2X7 U16934 ( .A(n4267), .B(n4278), .Z(n2981) );
  HS65_LL_NAND2X7 U16935 ( .A(n4325), .B(n4338), .Z(n2846) );
  HS65_LL_NAND2X7 U16936 ( .A(n4216), .B(n4214), .Z(n3112) );
  HS65_LL_NAND2X7 U16937 ( .A(n5741), .B(n5738), .Z(n4485) );
  HS65_LL_NAND2X7 U16938 ( .A(n7333), .B(n7330), .Z(n6078) );
  HS65_LL_NAND2X7 U16939 ( .A(n5738), .B(n5748), .Z(n4552) );
  HS65_LL_NAND2X7 U16940 ( .A(n7330), .B(n7340), .Z(n6145) );
  HS65_LL_NAND2X7 U16941 ( .A(n4217), .B(n4203), .Z(n2855) );
  HS65_LL_NAND2X7 U16942 ( .A(n8925), .B(n8908), .Z(n8057) );
  HS65_LL_NAND2X7 U16943 ( .A(n8984), .B(n8985), .Z(n8302) );
  HS65_LL_NOR2X6 U16944 ( .A(n337), .B(n338), .Z(n8918) );
  HS65_LL_NOR2X6 U16945 ( .A(n159), .B(n160), .Z(n4137) );
  HS65_LL_NOR2X6 U16946 ( .A(n379), .B(n380), .Z(n8988) );
  HS65_LL_NOR2X6 U16947 ( .A(n331), .B(n336), .Z(n8925) );
  HS65_LL_NOR2X6 U16948 ( .A(n425), .B(n424), .Z(n4329) );
  HS65_LL_NOR2X6 U16949 ( .A(n595), .B(n594), .Z(n9043) );
  HS65_LL_NOR2X6 U16950 ( .A(n115), .B(n114), .Z(n9101) );
  HS65_LL_NOR2X6 U16951 ( .A(n632), .B(n641), .Z(n4271) );
  HS65_LL_NOR2X6 U16952 ( .A(n204), .B(n205), .Z(n4202) );
  HS65_LL_NOR2X6 U16953 ( .A(n358), .B(n359), .Z(n8932) );
  HS65_LL_NOR2X6 U16954 ( .A(n402), .B(n403), .Z(n8987) );
  HS65_LL_NOR2X6 U16955 ( .A(n445), .B(n446), .Z(n4331) );
  HS65_LL_NOR2X6 U16956 ( .A(n227), .B(n228), .Z(n4215) );
  HS65_LL_NAND2X7 U16957 ( .A(n4266), .B(n4281), .Z(n2876) );
  HS65_LL_NAND2X7 U16958 ( .A(n5920), .B(n5930), .Z(n5616) );
  HS65_LL_NAND2X7 U16959 ( .A(n5861), .B(n5871), .Z(n5591) );
  HS65_LL_NAND2X7 U16960 ( .A(n7454), .B(n7466), .Z(n7183) );
  HS65_LL_NAND2X7 U16961 ( .A(n7512), .B(n7522), .Z(n7208) );
  HS65_LL_NAND2X7 U16962 ( .A(n7404), .B(n7405), .Z(n7164) );
  HS65_LL_NAND2X7 U16963 ( .A(n1841), .B(n1854), .Z(n1745) );
  HS65_LL_NAND2X7 U16964 ( .A(n5865), .B(n5875), .Z(n4727) );
  HS65_LL_NAND2X7 U16965 ( .A(n5924), .B(n5934), .Z(n4789) );
  HS65_LL_NAND2X7 U16966 ( .A(n7516), .B(n7526), .Z(n6382) );
  HS65_LL_NAND2X7 U16967 ( .A(n7459), .B(n7468), .Z(n6343) );
  HS65_LL_NAND2X7 U16968 ( .A(n7398), .B(n7399), .Z(n6236) );
  HS65_LL_NAND2X7 U16969 ( .A(n5806), .B(n5807), .Z(n4643) );
  HS65_LL_NAND2X7 U16970 ( .A(n4325), .B(n4343), .Z(n2829) );
  HS65_LL_NAND2X7 U16971 ( .A(n4216), .B(n4209), .Z(n3097) );
  HS65_LL_NAND2X7 U16972 ( .A(n2593), .B(n2606), .Z(n2497) );
  HS65_LL_NAND2X7 U16973 ( .A(n2217), .B(n2230), .Z(n2121) );
  HS65_LL_NAND2X7 U16974 ( .A(n1465), .B(n1478), .Z(n1369) );
  HS65_LL_NAND2X7 U16975 ( .A(n4267), .B(n4280), .Z(n3134) );
  HS65_LL_NAND2X7 U16976 ( .A(n8916), .B(n8932), .Z(n8313) );
  HS65_LL_NAND2X7 U16977 ( .A(n4159), .B(n4151), .Z(n3588) );
  HS65_LL_NAND2X7 U16978 ( .A(n9047), .B(n9019), .Z(n8132) );
  HS65_LL_NAND2X7 U16979 ( .A(n9105), .B(n9077), .Z(n8183) );
  HS65_LL_NAND2X7 U16980 ( .A(n2232), .B(n2218), .Z(n2069) );
  HS65_LL_NAND2X7 U16981 ( .A(n1480), .B(n1466), .Z(n1317) );
  HS65_LL_NAND2X7 U16982 ( .A(n4284), .B(n4264), .Z(n3343) );
  HS65_LL_NAND2X7 U16983 ( .A(n5872), .B(n5851), .Z(n5604) );
  HS65_LL_NAND2X7 U16984 ( .A(n5931), .B(n5910), .Z(n5629) );
  HS65_LL_NAND2X7 U16985 ( .A(n7456), .B(n7443), .Z(n7196) );
  HS65_LL_NAND2X7 U16986 ( .A(n7523), .B(n7502), .Z(n7221) );
  HS65_LL_NAND2X7 U16987 ( .A(n7400), .B(n7396), .Z(n7170) );
  HS65_LL_NAND2X7 U16988 ( .A(n5808), .B(n5804), .Z(n5578) );
  HS65_LL_NAND2X7 U16989 ( .A(n4323), .B(n4338), .Z(n3204) );
  HS65_LL_NAND2X7 U16990 ( .A(n8978), .B(n8968), .Z(n7966) );
  HS65_LL_NAND2X7 U16991 ( .A(n7337), .B(n7332), .Z(n7094) );
  HS65_LL_NAND2X7 U16992 ( .A(n5745), .B(n5740), .Z(n5502) );
  HS65_LL_NAND2X7 U16993 ( .A(n8916), .B(n8930), .Z(n8357) );
  HS65_LL_NAND2X7 U16994 ( .A(n5924), .B(n5936), .Z(n4494) );
  HS65_LL_NAND2X7 U16995 ( .A(n5865), .B(n5877), .Z(n4455) );
  HS65_LL_NAND2X7 U16996 ( .A(n7516), .B(n7528), .Z(n6087) );
  HS65_LL_NAND2X7 U16997 ( .A(n7459), .B(n7460), .Z(n6048) );
  HS65_LL_NAND2X7 U16998 ( .A(n7398), .B(n7395), .Z(n6219) );
  HS65_LL_NAND2X7 U16999 ( .A(n5806), .B(n5803), .Z(n4626) );
  HS65_LL_NAND2X7 U17000 ( .A(n7512), .B(n7525), .Z(n6581) );
  HS65_LL_NAND2X7 U17001 ( .A(n7454), .B(n7461), .Z(n6469) );
  HS65_LL_NAND2X7 U17002 ( .A(n5861), .B(n5874), .Z(n4876) );
  HS65_LL_NAND2X7 U17003 ( .A(n5920), .B(n5933), .Z(n4988) );
  HS65_LL_NAND2X7 U17004 ( .A(n7404), .B(n7401), .Z(n6455) );
  HS65_LL_NAND2X7 U17005 ( .A(n5812), .B(n5809), .Z(n4862) );
  HS65_LL_NAND2X7 U17006 ( .A(n2608), .B(n2594), .Z(n2445) );
  HS65_LL_NAND2X7 U17007 ( .A(n4146), .B(n4158), .Z(n3253) );
  HS65_LL_NAND2X7 U17008 ( .A(n1856), .B(n1842), .Z(n1693) );
  HS65_LL_NAND2X7 U17009 ( .A(n5746), .B(n5747), .Z(n4567) );
  HS65_LL_NAND2X7 U17010 ( .A(n7338), .B(n7339), .Z(n6160) );
  HS65_LL_NAND2X7 U17011 ( .A(n2228), .B(n2209), .Z(n2146) );
  HS65_LL_NAND2X7 U17012 ( .A(n5746), .B(n5742), .Z(n5514) );
  HS65_LL_NAND2X7 U17013 ( .A(n7338), .B(n7334), .Z(n7106) );
  HS65_LL_NAND2X7 U17014 ( .A(n4209), .B(n4213), .Z(n3115) );
  HS65_LL_NAND2X7 U17015 ( .A(n5929), .B(n5930), .Z(n4492) );
  HS65_LL_NAND2X7 U17016 ( .A(n5870), .B(n5871), .Z(n4453) );
  HS65_LL_NAND2X7 U17017 ( .A(n7521), .B(n7522), .Z(n6085) );
  HS65_LL_NAND2X7 U17018 ( .A(n5805), .B(n5813), .Z(n4850) );
  HS65_LL_NAND2X7 U17019 ( .A(n7397), .B(n7405), .Z(n6443) );
  HS65_LL_NAND2X7 U17020 ( .A(n7453), .B(n7466), .Z(n6046) );
  HS65_LL_NAND2X7 U17021 ( .A(n4148), .B(n4155), .Z(n3994) );
  HS65_LL_NAND2X7 U17022 ( .A(n8929), .B(n8908), .Z(n8034) );
  HS65_LL_NAND2X7 U17023 ( .A(n2586), .B(n2587), .Z(n2240) );
  HS65_LL_NAND2X7 U17024 ( .A(n1834), .B(n1835), .Z(n1488) );
  HS65_LL_NAND2X7 U17025 ( .A(n9085), .B(n9086), .Z(n8169) );
  HS65_LL_NAND2X7 U17026 ( .A(n9027), .B(n9028), .Z(n8146) );
  HS65_LL_NAND2X7 U17027 ( .A(n2210), .B(n2211), .Z(n1864) );
  HS65_LL_NAND2X7 U17028 ( .A(n1458), .B(n1459), .Z(n1112) );
  HS65_LL_NAND2X7 U17029 ( .A(n9107), .B(n9078), .Z(n7650) );
  HS65_LL_NAND2X7 U17030 ( .A(n9049), .B(n9020), .Z(n7630) );
  HS65_LL_NAND2X7 U17031 ( .A(n1852), .B(n1833), .Z(n1770) );
  HS65_LL_NAND2X7 U17032 ( .A(n2604), .B(n2585), .Z(n2522) );
  HS65_LL_NAND2X7 U17033 ( .A(n1476), .B(n1457), .Z(n1394) );
  HS65_LL_NAND2X7 U17034 ( .A(n8989), .B(n8990), .Z(n7960) );
  HS65_LL_NAND2X7 U17035 ( .A(n1840), .B(n1855), .Z(n1519) );
  HS65_LL_NAND2X7 U17036 ( .A(n2592), .B(n2607), .Z(n2271) );
  HS65_LL_NAND2X7 U17037 ( .A(n1464), .B(n1479), .Z(n1143) );
  HS65_LL_NAND2X7 U17038 ( .A(n2216), .B(n2231), .Z(n1895) );
  HS65_LL_NAND2X7 U17039 ( .A(n5934), .B(n5935), .Z(n4500) );
  HS65_LL_NAND2X7 U17040 ( .A(n5875), .B(n5876), .Z(n4461) );
  HS65_LL_NAND2X7 U17041 ( .A(n7526), .B(n7527), .Z(n6093) );
  HS65_LL_NAND2X7 U17042 ( .A(n5807), .B(n5814), .Z(n5496) );
  HS65_LL_NAND2X7 U17043 ( .A(n7399), .B(n7406), .Z(n7088) );
  HS65_LL_NAND2X7 U17044 ( .A(n7468), .B(n7469), .Z(n6054) );
  HS65_LL_NAND2X7 U17045 ( .A(n9048), .B(n9046), .Z(n7836) );
  HS65_LL_NAND2X7 U17046 ( .A(n9106), .B(n9104), .Z(n7875) );
  HS65_LL_NAND2X7 U17047 ( .A(n5744), .B(n5741), .Z(n4550) );
  HS65_LL_NAND2X7 U17048 ( .A(n7336), .B(n7333), .Z(n6143) );
  HS65_LL_NAND2X7 U17049 ( .A(n9042), .B(n9041), .Z(n7631) );
  HS65_LL_NAND2X7 U17050 ( .A(n9100), .B(n9099), .Z(n7651) );
  HS65_LL_NAND2X7 U17051 ( .A(n4217), .B(n4212), .Z(n2956) );
  HS65_LL_NAND2X7 U17052 ( .A(n5913), .B(n5923), .Z(n4775) );
  HS65_LL_NAND2X7 U17053 ( .A(n7505), .B(n7515), .Z(n6368) );
  HS65_LL_NAND2X7 U17054 ( .A(n5854), .B(n5864), .Z(n4733) );
  HS65_LL_NAND2X7 U17055 ( .A(n7446), .B(n7458), .Z(n6329) );
  HS65_LL_NAND2X7 U17056 ( .A(n7392), .B(n7402), .Z(n6222) );
  HS65_LL_NAND2X7 U17057 ( .A(n5800), .B(n5810), .Z(n4629) );
  HS65_LL_NAND2X7 U17058 ( .A(n9102), .B(n9109), .Z(n7919) );
  HS65_LL_NAND2X7 U17059 ( .A(n9044), .B(n9051), .Z(n7821) );
  HS65_LL_NAND2X7 U17060 ( .A(n5864), .B(n5876), .Z(n4593) );
  HS65_LL_NAND2X7 U17061 ( .A(n5923), .B(n5935), .Z(n4610) );
  HS65_LL_NAND2X7 U17062 ( .A(n7515), .B(n7527), .Z(n6203) );
  HS65_LL_NAND2X7 U17063 ( .A(n7458), .B(n7469), .Z(n6186) );
  HS65_LL_NAND2X7 U17064 ( .A(n5742), .B(n5728), .Z(n4668) );
  HS65_LL_NAND2X7 U17065 ( .A(n7334), .B(n7320), .Z(n6261) );
  HS65_LL_NAND2X7 U17066 ( .A(n7503), .B(n7522), .Z(n6094) );
  HS65_LL_NAND2X7 U17067 ( .A(n7444), .B(n7466), .Z(n6055) );
  HS65_LL_NAND2X7 U17068 ( .A(n5852), .B(n5871), .Z(n4462) );
  HS65_LL_NAND2X7 U17069 ( .A(n5911), .B(n5930), .Z(n4501) );
  HS65_LL_NAND2X7 U17070 ( .A(n5790), .B(n5813), .Z(n4523) );
  HS65_LL_NAND2X7 U17071 ( .A(n5728), .B(n5751), .Z(n4483) );
  HS65_LL_NAND2X7 U17072 ( .A(n7382), .B(n7405), .Z(n6116) );
  HS65_LL_NAND2X7 U17073 ( .A(n7320), .B(n7343), .Z(n6076) );
  HS65_LL_NAND2X7 U17074 ( .A(n4328), .B(n4327), .Z(n2993) );
  HS65_LL_NAND2X7 U17075 ( .A(n4269), .B(n4268), .Z(n2968) );
  HS65_LL_NAND2X7 U17076 ( .A(n4147), .B(n4158), .Z(n3224) );
  HS65_LL_NAND2X7 U17077 ( .A(n4213), .B(n4214), .Z(n2939) );
  HS65_LL_NAND2X7 U17078 ( .A(n5931), .B(n5930), .Z(n4508) );
  HS65_LL_NAND2X7 U17079 ( .A(n5872), .B(n5871), .Z(n4447) );
  HS65_LL_NAND2X7 U17080 ( .A(n7523), .B(n7522), .Z(n6101) );
  HS65_LL_NAND2X7 U17081 ( .A(n5808), .B(n5813), .Z(n4654) );
  HS65_LL_NAND2X7 U17082 ( .A(n7400), .B(n7405), .Z(n6247) );
  HS65_LL_NAND2X7 U17083 ( .A(n7456), .B(n7466), .Z(n6040) );
  HS65_LL_NAND2X7 U17084 ( .A(n2206), .B(n2232), .Z(n1861) );
  HS65_LL_NAND2X7 U17085 ( .A(n1464), .B(n1474), .Z(n1162) );
  HS65_LL_NAND2X7 U17086 ( .A(n2216), .B(n2226), .Z(n1914) );
  HS65_LL_NAND2X7 U17087 ( .A(n1454), .B(n1480), .Z(n1109) );
  HS65_LL_NAND2X7 U17088 ( .A(n1830), .B(n1856), .Z(n1485) );
  HS65_LL_NAND2X7 U17089 ( .A(n2582), .B(n2608), .Z(n2237) );
  HS65_LL_NAND2X7 U17090 ( .A(n4326), .B(n4337), .Z(n3184) );
  HS65_LL_NAND2X7 U17091 ( .A(n5727), .B(n5728), .Z(n4549) );
  HS65_LL_NAND2X7 U17092 ( .A(n7319), .B(n7320), .Z(n6142) );
  HS65_LL_NAND2X7 U17093 ( .A(n4145), .B(n4146), .Z(n3048) );
  HS65_LL_NAND2X7 U17094 ( .A(n4154), .B(n4152), .Z(n3042) );
  HS65_LL_NAND2X7 U17095 ( .A(n4266), .B(n4272), .Z(n2890) );
  HS65_LL_NAND2X7 U17096 ( .A(n8931), .B(n8911), .Z(n7940) );
  HS65_LL_NAND2X7 U17097 ( .A(n4269), .B(n4270), .Z(n2884) );
  HS65_LL_NAND2X7 U17098 ( .A(n5750), .B(n5751), .Z(n5508) );
  HS65_LL_NAND2X7 U17099 ( .A(n7342), .B(n7343), .Z(n7100) );
  HS65_LL_NAND2X7 U17100 ( .A(n9103), .B(n9104), .Z(n7653) );
  HS65_LL_NAND2X7 U17101 ( .A(n9045), .B(n9046), .Z(n7633) );
  HS65_LL_NAND2X7 U17102 ( .A(n9040), .B(n9028), .Z(n7622) );
  HS65_LL_NAND2X7 U17103 ( .A(n9098), .B(n9086), .Z(n7662) );
  HS65_LL_NAND2X7 U17104 ( .A(n1840), .B(n1850), .Z(n1538) );
  HS65_LL_NAND2X7 U17105 ( .A(n2592), .B(n2602), .Z(n2290) );
  HS65_LL_NAND2X7 U17106 ( .A(n8916), .B(n8917), .Z(n8527) );
  HS65_LL_NAND2X7 U17107 ( .A(n4266), .B(n4284), .Z(n2881) );
  HS65_LL_NAND2X7 U17108 ( .A(n1834), .B(n1841), .Z(n1520) );
  HS65_LL_NAND2X7 U17109 ( .A(n2586), .B(n2593), .Z(n2272) );
  HS65_LL_NAND2X7 U17110 ( .A(n1458), .B(n1465), .Z(n1144) );
  HS65_LL_NAND2X7 U17111 ( .A(n2210), .B(n2217), .Z(n1896) );
  HS65_LL_NAND2X7 U17112 ( .A(n8984), .B(n8987), .Z(n8067) );
  HS65_LL_NAND2X7 U17113 ( .A(n4158), .B(n4155), .Z(n3054) );
  HS65_LL_NOR2X6 U17114 ( .A(n917), .B(n918), .Z(n2587) );
  HS65_LL_NOR2X6 U17115 ( .A(n835), .B(n836), .Z(n1835) );
  HS65_LL_NAND2X7 U17116 ( .A(n4211), .B(n4201), .Z(n2932) );
  HS65_LL_NAND2X7 U17117 ( .A(n1835), .B(n1854), .Z(n1532) );
  HS65_LL_NOR2X6 U17118 ( .A(n794), .B(n795), .Z(n2211) );
  HS65_LL_NOR2X6 U17119 ( .A(n876), .B(n877), .Z(n1459) );
  HS65_LL_NAND2X7 U17120 ( .A(n4329), .B(n4341), .Z(n3192) );
  HS65_LL_NAND2X7 U17121 ( .A(n4212), .B(n4220), .Z(n2926) );
  HS65_LL_NAND2X7 U17122 ( .A(n2604), .B(n2603), .Z(n2520) );
  HS65_LL_NAND2X7 U17123 ( .A(n2587), .B(n2606), .Z(n2284) );
  HS65_LL_NAND2X7 U17124 ( .A(n2211), .B(n2230), .Z(n1908) );
  HS65_LL_NAND2X7 U17125 ( .A(n1459), .B(n1478), .Z(n1156) );
  HS65_LL_NAND2X7 U17126 ( .A(n2228), .B(n2227), .Z(n2144) );
  HS65_LL_NAND2X7 U17127 ( .A(n1476), .B(n1475), .Z(n1392) );
  HS65_LL_NAND2X7 U17128 ( .A(n4343), .B(n4323), .Z(n3397) );
  HS65_LL_NAND2X7 U17129 ( .A(n1852), .B(n1851), .Z(n1768) );
  HS65_LL_NAND2X7 U17130 ( .A(n4339), .B(n4324), .Z(n3972) );
  HS65_LL_NAND2X7 U17131 ( .A(n9027), .B(n9041), .Z(n7807) );
  HS65_LL_NAND2X7 U17132 ( .A(n9085), .B(n9099), .Z(n7905) );
  HS65_LL_NAND2X7 U17133 ( .A(n5743), .B(n5751), .Z(n4712) );
  HS65_LL_NAND2X7 U17134 ( .A(n7335), .B(n7343), .Z(n6305) );
  HS65_LL_NAND2X7 U17135 ( .A(n4340), .B(n4338), .Z(n3193) );
  HS65_LL_NAND2X7 U17136 ( .A(n4221), .B(n4214), .Z(n2927) );
  HS65_LL_NAND2X7 U17137 ( .A(n4270), .B(n4277), .Z(n3128) );
  HS65_LL_NAND2X7 U17138 ( .A(n4210), .B(n4214), .Z(n3926) );
  HS65_LL_NAND2X7 U17139 ( .A(n4339), .B(n4338), .Z(n3970) );
  HS65_LL_NAND2X7 U17140 ( .A(n8918), .B(n8919), .Z(n8028) );
  HS65_LL_NAND2X7 U17141 ( .A(n2229), .B(n2227), .Z(n1909) );
  HS65_LL_NAND2X7 U17142 ( .A(n1477), .B(n1475), .Z(n1157) );
  HS65_LL_NAND2X7 U17143 ( .A(n9040), .B(n9048), .Z(n8421) );
  HS65_LL_NAND2X7 U17144 ( .A(n9098), .B(n9106), .Z(n8473) );
  HS65_LL_NOR2X6 U17145 ( .A(n381), .B(n382), .Z(n8989) );
  HS65_LL_NAND2X7 U17146 ( .A(n2594), .B(n2603), .Z(n2297) );
  HS65_LL_NAND2X7 U17147 ( .A(n4282), .B(n4265), .Z(n3952) );
  HS65_LL_NAND2X7 U17148 ( .A(n2218), .B(n2227), .Z(n1921) );
  HS65_LL_NAND2X7 U17149 ( .A(n1466), .B(n1475), .Z(n1169) );
  HS65_LL_NAND2X7 U17150 ( .A(n2605), .B(n2603), .Z(n2285) );
  HS65_LL_NAND2X7 U17151 ( .A(n8986), .B(n8971), .Z(n7858) );
  HS65_LL_NOR2X6 U17152 ( .A(n116), .B(n117), .Z(n9078) );
  HS65_LL_NOR2X6 U17153 ( .A(n596), .B(n597), .Z(n9020) );
  HS65_LL_NAND2X7 U17154 ( .A(n4282), .B(n4281), .Z(n3950) );
  HS65_LL_NAND2X7 U17155 ( .A(n4283), .B(n4281), .Z(n3129) );
  HS65_LL_NAND2X7 U17156 ( .A(n4210), .B(n4219), .Z(n3928) );
  HS65_LL_NAND2X7 U17157 ( .A(n1853), .B(n1851), .Z(n1533) );
  HS65_LL_NAND2X7 U17158 ( .A(n5748), .B(n5752), .Z(n5013) );
  HS65_LL_NAND2X7 U17159 ( .A(n7340), .B(n7344), .Z(n6606) );
  HS65_LL_NAND2X7 U17160 ( .A(n9019), .B(n9020), .Z(n8128) );
  HS65_LL_NAND2X7 U17161 ( .A(n9077), .B(n9078), .Z(n8179) );
  HS65_LL_NAND2X7 U17162 ( .A(n1842), .B(n1851), .Z(n1545) );
  HS65_LL_NAND2X7 U17163 ( .A(n5746), .B(n5751), .Z(n4685) );
  HS65_LL_NAND2X7 U17164 ( .A(n7338), .B(n7343), .Z(n6278) );
  HS65_LL_NAND2X7 U17165 ( .A(n8970), .B(n8991), .Z(n7961) );
  HS65_LL_NAND2X7 U17166 ( .A(n8910), .B(n8930), .Z(n8029) );
  HS65_LL_NAND2X7 U17167 ( .A(n5875), .B(n5854), .Z(n4732) );
  HS65_LL_NAND2X7 U17168 ( .A(n5934), .B(n5913), .Z(n4794) );
  HS65_LL_NAND2X7 U17169 ( .A(n7526), .B(n7505), .Z(n6387) );
  HS65_LL_NAND2X7 U17170 ( .A(n7468), .B(n7446), .Z(n6348) );
  HS65_LL_NAND2X7 U17171 ( .A(n7399), .B(n7392), .Z(n6241) );
  HS65_LL_NAND2X7 U17172 ( .A(n5807), .B(n5800), .Z(n4648) );
  HS65_LL_NAND2X7 U17173 ( .A(n5872), .B(n5874), .Z(n4728) );
  HS65_LL_NAND2X7 U17174 ( .A(n5931), .B(n5933), .Z(n4790) );
  HS65_LL_NAND2X7 U17175 ( .A(n7523), .B(n7525), .Z(n6383) );
  HS65_LL_NAND2X7 U17176 ( .A(n7456), .B(n7461), .Z(n6344) );
  HS65_LL_NAND2X7 U17177 ( .A(n7400), .B(n7401), .Z(n6237) );
  HS65_LL_NAND2X7 U17178 ( .A(n5808), .B(n5809), .Z(n4644) );
  HS65_LL_NAND2X7 U17179 ( .A(n9103), .B(n9098), .Z(n8018) );
  HS65_LL_NAND2X7 U17180 ( .A(n5745), .B(n5738), .Z(n4571) );
  HS65_LL_NAND2X7 U17181 ( .A(n7337), .B(n7330), .Z(n6164) );
  HS65_LL_NAND2X7 U17182 ( .A(n5920), .B(n5910), .Z(n4608) );
  HS65_LL_NAND2X7 U17183 ( .A(n5861), .B(n5851), .Z(n4591) );
  HS65_LL_NAND2X7 U17184 ( .A(n5812), .B(n5804), .Z(n4524) );
  HS65_LL_NAND2X7 U17185 ( .A(n7512), .B(n7502), .Z(n6201) );
  HS65_LL_NAND2X7 U17186 ( .A(n7404), .B(n7396), .Z(n6117) );
  HS65_LL_NAND2X7 U17187 ( .A(n7454), .B(n7443), .Z(n6184) );
  HS65_LL_NAND2X7 U17188 ( .A(n9099), .B(n9104), .Z(n7882) );
  HS65_LL_NAND2X7 U17189 ( .A(n9041), .B(n9046), .Z(n7783) );
  HS65_LL_NAND2X7 U17190 ( .A(n4209), .B(n4210), .Z(n2933) );
  HS65_LL_NAND2X7 U17191 ( .A(n2207), .B(n2229), .Z(n1920) );
  HS65_LL_NAND2X7 U17192 ( .A(n1455), .B(n1477), .Z(n1168) );
  HS65_LL_NOR2X6 U17193 ( .A(n900), .B(n899), .Z(n2582) );
  HS65_LL_NOR2X6 U17194 ( .A(n818), .B(n817), .Z(n1830) );
  HS65_LL_NOR2X6 U17195 ( .A(n859), .B(n858), .Z(n1454) );
  HS65_LL_NOR2X6 U17196 ( .A(n777), .B(n776), .Z(n2206) );
  HS65_LL_NAND2X7 U17197 ( .A(n2583), .B(n2605), .Z(n2296) );
  HS65_LL_NAND2X7 U17198 ( .A(n1831), .B(n1853), .Z(n1544) );
  HS65_LL_NAND2X7 U17199 ( .A(n5742), .B(n5743), .Z(n4572) );
  HS65_LL_NAND2X7 U17200 ( .A(n7334), .B(n7335), .Z(n6165) );
  HS65_LL_NAND2X7 U17201 ( .A(n2608), .B(n2604), .Z(n2291) );
  HS65_LL_NAND2X7 U17202 ( .A(n2232), .B(n2228), .Z(n1915) );
  HS65_LL_NAND2X7 U17203 ( .A(n1480), .B(n1476), .Z(n1163) );
  HS65_LL_NAND2X7 U17204 ( .A(n1834), .B(n1855), .Z(n1505) );
  HS65_LL_NAND2X7 U17205 ( .A(n2586), .B(n2607), .Z(n2257) );
  HS65_LL_NAND2X7 U17206 ( .A(n1458), .B(n1479), .Z(n1129) );
  HS65_LL_NAND2X7 U17207 ( .A(n2210), .B(n2231), .Z(n1881) );
  HS65_LL_NAND2X7 U17208 ( .A(n1841), .B(n1844), .Z(n1521) );
  HS65_LL_NAND2X7 U17209 ( .A(n2593), .B(n2596), .Z(n2273) );
  HS65_LL_NAND2X7 U17210 ( .A(n1465), .B(n1468), .Z(n1145) );
  HS65_LL_NAND2X7 U17211 ( .A(n2217), .B(n2220), .Z(n1897) );
  HS65_LL_NAND2X7 U17212 ( .A(n4327), .B(n4330), .Z(n2994) );
  HS65_LL_NAND2X7 U17213 ( .A(n1856), .B(n1852), .Z(n1539) );
  HS65_LL_NAND2X7 U17214 ( .A(n4215), .B(n4221), .Z(n2938) );
  HS65_LL_NAND2X7 U17215 ( .A(n4331), .B(n4340), .Z(n3203) );
  HS65_LL_NOR2X6 U17216 ( .A(n662), .B(n663), .Z(n4266) );
  HS65_LL_NAND2X7 U17217 ( .A(n8932), .B(n8910), .Z(n7942) );
  HS65_LL_NOR2X6 U17218 ( .A(n643), .B(n642), .Z(n4270) );
  HS65_LL_NOR2X6 U17219 ( .A(n207), .B(n206), .Z(n4212) );
  HS65_LL_NAND2X7 U17220 ( .A(n4284), .B(n4282), .Z(n3135) );
  HS65_LL_NAND2X7 U17221 ( .A(n4328), .B(n4342), .Z(n2845) );
  HS65_LL_NAND2X7 U17222 ( .A(n4269), .B(n4278), .Z(n2875) );
  HS65_LL_NAND2X7 U17223 ( .A(n8987), .B(n8970), .Z(n7860) );
  HS65_LL_NAND2X7 U17224 ( .A(n5910), .B(n5929), .Z(n4795) );
  HS65_LL_NAND2X7 U17225 ( .A(n5851), .B(n5870), .Z(n4734) );
  HS65_LL_NAND2X7 U17226 ( .A(n5804), .B(n5805), .Z(n4649) );
  HS65_LL_NAND2X7 U17227 ( .A(n7502), .B(n7521), .Z(n6388) );
  HS65_LL_NAND2X7 U17228 ( .A(n7396), .B(n7397), .Z(n6242) );
  HS65_LL_NAND2X7 U17229 ( .A(n7443), .B(n7453), .Z(n6349) );
  HS65_LL_NAND2X7 U17230 ( .A(n2607), .B(n2596), .Z(n2333) );
  HS65_LL_NAND2X7 U17231 ( .A(n1855), .B(n1844), .Z(n1581) );
  HS65_LL_NAND2X7 U17232 ( .A(n8988), .B(n8979), .Z(n7847) );
  HS65_LL_NAND2X7 U17233 ( .A(n2231), .B(n2220), .Z(n1957) );
  HS65_LL_NAND2X7 U17234 ( .A(n1479), .B(n1468), .Z(n1205) );
  HS65_LL_NAND2X7 U17235 ( .A(n2218), .B(n2209), .Z(n1863) );
  HS65_LL_NAND2X7 U17236 ( .A(n8928), .B(n8907), .Z(n7767) );
  HS65_LL_NOR2X6 U17237 ( .A(n161), .B(n162), .Z(n4152) );
  HS65_LL_NOR2X6 U17238 ( .A(n133), .B(n138), .Z(n9104) );
  HS65_LL_NOR2X6 U17239 ( .A(n613), .B(n618), .Z(n9046) );
  HS65_LL_NAND2X7 U17240 ( .A(n1842), .B(n1833), .Z(n1487) );
  HS65_LL_NAND2X7 U17241 ( .A(n2594), .B(n2585), .Z(n2239) );
  HS65_LL_NAND2X7 U17242 ( .A(n1466), .B(n1457), .Z(n1111) );
  HS65_LL_NAND2X7 U17243 ( .A(n4203), .B(n4202), .Z(n2856) );
  HS65_LL_NAND2X7 U17244 ( .A(n4268), .B(n4271), .Z(n2969) );
  HS65_LL_NAND2X7 U17245 ( .A(n4217), .B(n4218), .Z(n2940) );
  HS65_LL_NAND2X7 U17246 ( .A(n8925), .B(n8926), .Z(n7948) );
  HS65_LL_NAND2X7 U17247 ( .A(n4323), .B(n4324), .Z(n2831) );
  HS65_LL_NAND2X7 U17248 ( .A(n8977), .B(n8967), .Z(n7749) );
  HS65_LL_NAND2X7 U17249 ( .A(n4218), .B(n4202), .Z(n3067) );
  HS65_LL_NAND2X7 U17250 ( .A(n4343), .B(n4339), .Z(n3198) );
  HS65_LL_NAND2X7 U17251 ( .A(n4342), .B(n4330), .Z(n3412) );
  HS65_LL_NAND2X7 U17252 ( .A(n5750), .B(n5742), .Z(n4484) );
  HS65_LL_NAND2X7 U17253 ( .A(n7342), .B(n7334), .Z(n6077) );
  HS65_LL_NAND2X7 U17254 ( .A(n2209), .B(n2229), .Z(n1951) );
  HS65_LL_NAND2X7 U17255 ( .A(n1457), .B(n1477), .Z(n1199) );
  HS65_LL_NAND2X7 U17256 ( .A(n8926), .B(n8907), .Z(n7947) );
  HS65_LL_NAND2X7 U17257 ( .A(n4272), .B(n4264), .Z(n3157) );
  HS65_LL_NAND2X7 U17258 ( .A(n4272), .B(n4283), .Z(n3140) );
  HS65_LL_NAND2X7 U17259 ( .A(n1480), .B(n1477), .Z(n1180) );
  HS65_LL_NAND2X7 U17260 ( .A(n2232), .B(n2229), .Z(n1932) );
  HS65_LL_NAND2X7 U17261 ( .A(n8931), .B(n8930), .Z(n8630) );
  HS65_LL_NAND2X7 U17262 ( .A(n8986), .B(n8991), .Z(n8649) );
  HS65_LL_NAND2X7 U17263 ( .A(n8916), .B(n8911), .Z(n7769) );
  HS65_LL_NAND2X7 U17264 ( .A(n9043), .B(n9047), .Z(n8155) );
  HS65_LL_NAND2X7 U17265 ( .A(n9101), .B(n9105), .Z(n8178) );
  HS65_LL_NAND2X7 U17266 ( .A(n4264), .B(n4265), .Z(n2883) );
  HS65_LL_NAND2X7 U17267 ( .A(n2585), .B(n2605), .Z(n2327) );
  HS65_LL_NAND2X7 U17268 ( .A(n1850), .B(n1844), .Z(n1609) );
  HS65_LL_NAND2X7 U17269 ( .A(n2602), .B(n2596), .Z(n2361) );
  HS65_LL_NAND2X7 U17270 ( .A(n2226), .B(n2220), .Z(n1985) );
  HS65_LL_NAND2X7 U17271 ( .A(n1474), .B(n1468), .Z(n1233) );
  HS65_LL_NAND2X7 U17272 ( .A(n4326), .B(n4327), .Z(n2997) );
  HS65_LL_NAND2X7 U17273 ( .A(n4267), .B(n4268), .Z(n2972) );
  HS65_LL_NAND2X7 U17274 ( .A(n4211), .B(n4203), .Z(n2859) );
  HS65_LL_NAND2X7 U17275 ( .A(n9101), .B(n9102), .Z(n8173) );
  HS65_LL_NAND2X7 U17276 ( .A(n9043), .B(n9044), .Z(n8150) );
  HS65_LL_NAND2X7 U17277 ( .A(n9102), .B(n9107), .Z(n7713) );
  HS65_LL_NAND2X7 U17278 ( .A(n9044), .B(n9049), .Z(n7675) );
  HS65_LL_NAND2X7 U17279 ( .A(n4201), .B(n4202), .Z(n3096) );
  HS65_LL_NAND2X7 U17280 ( .A(n4213), .B(n4219), .Z(n3095) );
  HS65_LL_NAND2X7 U17281 ( .A(n2608), .B(n2605), .Z(n2308) );
  HS65_LL_NAND2X7 U17282 ( .A(n8918), .B(n8907), .Z(n7943) );
  HS65_LL_NAND2X7 U17283 ( .A(n4337), .B(n4330), .Z(n3380) );
  HS65_LL_NAND2X7 U17284 ( .A(n8919), .B(n8928), .Z(n7941) );
  HS65_LL_NAND2X7 U17285 ( .A(n8988), .B(n8977), .Z(n8123) );
  HS65_LL_NAND2X7 U17286 ( .A(n8925), .B(n8928), .Z(n8369) );
  HS65_LL_NAND2X7 U17287 ( .A(n1833), .B(n1853), .Z(n1575) );
  HS65_LL_NAND2X7 U17288 ( .A(n4269), .B(n4280), .Z(n2888) );
  HS65_LL_NAND2X7 U17289 ( .A(n9034), .B(n9051), .Z(n7686) );
  HS65_LL_NAND2X7 U17290 ( .A(n9092), .B(n9109), .Z(n7724) );
  HS65_LL_NAND2X7 U17291 ( .A(n9045), .B(n9042), .Z(n7831) );
  HS65_LL_NAND2X7 U17292 ( .A(n8979), .B(n8967), .Z(n7846) );
  HS65_LL_NAND2X7 U17293 ( .A(n4324), .B(n4340), .Z(n3406) );
  HS65_LL_NAND2X7 U17294 ( .A(n5920), .B(n5921), .Z(n4495) );
  HS65_LL_NAND2X7 U17295 ( .A(n5861), .B(n5862), .Z(n4456) );
  HS65_LL_NAND2X7 U17296 ( .A(n7512), .B(n7513), .Z(n6088) );
  HS65_LL_NAND2X7 U17297 ( .A(n7454), .B(n7455), .Z(n6049) );
  HS65_LL_NAND2X7 U17298 ( .A(n4328), .B(n4337), .Z(n2836) );
  HS65_LL_NAND2X7 U17299 ( .A(n1856), .B(n1853), .Z(n1556) );
  HS65_LL_NAND2X7 U17300 ( .A(n8987), .B(n8992), .Z(n7980) );
  HS65_LL_NAND2X7 U17301 ( .A(n8932), .B(n8924), .Z(n8048) );
  HS65_LL_NAND2X7 U17302 ( .A(n8930), .B(n8924), .Z(n8039) );
  HS65_LL_NAND2X7 U17303 ( .A(n8929), .B(n8928), .Z(n8510) );
  HS65_LL_NAND2X7 U17304 ( .A(n8991), .B(n8992), .Z(n7971) );
  HS65_LL_NAND2X7 U17305 ( .A(n4209), .B(n4221), .Z(n2958) );
  HS65_LL_NAND2X7 U17306 ( .A(n4343), .B(n4340), .Z(n3185) );
  HS65_LL_NAND2X7 U17307 ( .A(n2206), .B(n2209), .Z(n2119) );
  HS65_LL_NAND2X7 U17308 ( .A(n5741), .B(n5752), .Z(n4670) );
  HS65_LL_NAND2X7 U17309 ( .A(n7333), .B(n7344), .Z(n6263) );
  HS65_LL_NAND2X7 U17310 ( .A(n8926), .B(n8919), .Z(n7768) );
  HS65_LL_NAND2X7 U17311 ( .A(n4341), .B(n4342), .Z(n2837) );
  HS65_LL_NAND2X7 U17312 ( .A(n4220), .B(n4218), .Z(n3116) );
  HS65_LL_NAND2X7 U17313 ( .A(n4277), .B(n4278), .Z(n2889) );
  HS65_LL_NAND2X7 U17314 ( .A(n2582), .B(n2585), .Z(n2495) );
  HS65_LL_NAND2X7 U17315 ( .A(n1454), .B(n1457), .Z(n1367) );
  HS65_LL_NAND2X7 U17316 ( .A(n1830), .B(n1833), .Z(n1743) );
  HS65_LL_NAND2X7 U17317 ( .A(n8978), .B(n8989), .Z(n8254) );
  HS65_LL_NAND2X7 U17318 ( .A(n4325), .B(n4324), .Z(n3807) );
  HS65_LL_NAND2X7 U17319 ( .A(n8929), .B(n8918), .Z(n8556) );
  HS65_LL_NAND2X7 U17320 ( .A(n8985), .B(n8992), .Z(n8106) );
  HS65_LL_NAND2X7 U17321 ( .A(n1850), .B(n1854), .Z(n1537) );
  HS65_LL_NAND2X7 U17322 ( .A(n8978), .B(n8977), .Z(n8207) );
  HS65_LL_NAND2X7 U17323 ( .A(n4326), .B(n4329), .Z(n3846) );
  HS65_LL_NAND2X7 U17324 ( .A(n2606), .B(n2607), .Z(n2245) );
  HS65_LL_NAND2X7 U17325 ( .A(n1854), .B(n1855), .Z(n1493) );
  HS65_LL_NAND2X7 U17326 ( .A(n1478), .B(n1479), .Z(n1117) );
  HS65_LL_NAND2X7 U17327 ( .A(n2230), .B(n2231), .Z(n1869) );
  HS65_LL_NAND2X7 U17328 ( .A(n4337), .B(n4341), .Z(n3197) );
  HS65_LL_NAND2X7 U17329 ( .A(n4201), .B(n4220), .Z(n2931) );
  HS65_LL_NAND2X7 U17330 ( .A(n9078), .B(n9109), .Z(n8776) );
  HS65_LL_NAND2X7 U17331 ( .A(n9020), .B(n9051), .Z(n8686) );
  HS65_LL_NAND2X7 U17332 ( .A(n9047), .B(n9051), .Z(n7624) );
  HS65_LL_NAND2X7 U17333 ( .A(n9105), .B(n9109), .Z(n7664) );
  HS65_LL_NAND2X7 U17334 ( .A(n5936), .B(n5913), .Z(n4499) );
  HS65_LL_NAND2X7 U17335 ( .A(n7528), .B(n7505), .Z(n6092) );
  HS65_LL_NAND2X7 U17336 ( .A(n5877), .B(n5854), .Z(n4460) );
  HS65_LL_NAND2X7 U17337 ( .A(n7460), .B(n7446), .Z(n6053) );
  HS65_LL_NAND2X7 U17338 ( .A(n5746), .B(n5727), .Z(n5507) );
  HS65_LL_NAND2X7 U17339 ( .A(n7338), .B(n7319), .Z(n7099) );
  HS65_LL_NAND2X7 U17340 ( .A(n8990), .B(n8977), .Z(n7859) );
  HS65_LL_NAND2X7 U17341 ( .A(n7339), .B(n7320), .Z(n7093) );
  HS65_LL_NAND2X7 U17342 ( .A(n5747), .B(n5728), .Z(n5501) );
  HS65_LL_NAND2X7 U17343 ( .A(n4219), .B(n4221), .Z(n3061) );
  HS65_LL_NAND2X7 U17344 ( .A(n2602), .B(n2606), .Z(n2289) );
  HS65_LL_NAND2X7 U17345 ( .A(n8967), .B(n8968), .Z(n8238) );
  HS65_LL_NAND2X7 U17346 ( .A(n5931), .B(n5921), .Z(n5555) );
  HS65_LL_NAND2X7 U17347 ( .A(n7523), .B(n7513), .Z(n7147) );
  HS65_LL_NAND2X7 U17348 ( .A(n5872), .B(n5862), .Z(n5533) );
  HS65_LL_NAND2X7 U17349 ( .A(n7456), .B(n7455), .Z(n7125) );
  HS65_LL_NAND2X7 U17350 ( .A(n5808), .B(n5789), .Z(n5571) );
  HS65_LL_NAND2X7 U17351 ( .A(n7400), .B(n7381), .Z(n7163) );
  HS65_LL_NAND2X7 U17352 ( .A(n4278), .B(n4271), .Z(n3299) );
  HS65_LL_NAND2X7 U17353 ( .A(n8911), .B(n8924), .Z(n8058) );
  HS65_LL_NAND2X7 U17354 ( .A(n2226), .B(n2230), .Z(n1913) );
  HS65_LL_NAND2X7 U17355 ( .A(n1474), .B(n1478), .Z(n1161) );
  HS65_LL_NAND2X7 U17356 ( .A(n4215), .B(n4213), .Z(n2957) );
  HS65_LL_NAND2X7 U17357 ( .A(n4331), .B(n4323), .Z(n3183) );
  HS65_LL_NAND2X7 U17358 ( .A(n4284), .B(n4283), .Z(n3158) );
  HS65_LL_NAND2X7 U17359 ( .A(n8985), .B(n8970), .Z(n8117) );
  HS65_LL_NAND2X7 U17360 ( .A(n8917), .B(n8910), .Z(n8363) );
  HS65_LL_NAND2X7 U17361 ( .A(n1455), .B(n1466), .Z(n1179) );
  HS65_LL_NAND2X7 U17362 ( .A(n2207), .B(n2218), .Z(n1931) );
  HS65_LL_NAND2X7 U17363 ( .A(n5936), .B(n5935), .Z(n4509) );
  HS65_LL_NAND2X7 U17364 ( .A(n7528), .B(n7527), .Z(n6102) );
  HS65_LL_NAND2X7 U17365 ( .A(n5877), .B(n5876), .Z(n4448) );
  HS65_LL_NAND2X7 U17366 ( .A(n7460), .B(n7469), .Z(n6041) );
  HS65_LL_NAND2X7 U17367 ( .A(n9040), .B(n9041), .Z(n7623) );
  HS65_LL_NAND2X7 U17368 ( .A(n9098), .B(n9099), .Z(n7663) );
  HS65_LL_NAND2X7 U17369 ( .A(n5922), .B(n5914), .Z(n4975) );
  HS65_LL_NAND2X7 U17370 ( .A(n5863), .B(n5855), .Z(n4922) );
  HS65_LL_NAND2X7 U17371 ( .A(n7514), .B(n7506), .Z(n6568) );
  HS65_LL_NAND2X7 U17372 ( .A(n7457), .B(n7447), .Z(n6515) );
  HS65_LL_NAND2X7 U17373 ( .A(n4268), .B(n4277), .Z(n3342) );
  HS65_LL_NAND2X7 U17374 ( .A(n1840), .B(n1835), .Z(n1695) );
  HS65_LL_NAND2X7 U17375 ( .A(n2592), .B(n2587), .Z(n2447) );
  HS65_LL_NAND2X7 U17376 ( .A(n1464), .B(n1459), .Z(n1319) );
  HS65_LL_NAND2X7 U17377 ( .A(n2216), .B(n2211), .Z(n2071) );
  HS65_LL_NAND2X7 U17378 ( .A(n8931), .B(n8932), .Z(n7949) );
  HS65_LL_NAND2X7 U17379 ( .A(n8910), .B(n8911), .Z(n8049) );
  HS65_LL_NAND2X7 U17380 ( .A(n2583), .B(n2594), .Z(n2307) );
  HS65_LL_NAND2X7 U17381 ( .A(n4327), .B(n4341), .Z(n3396) );
  HS65_LL_NAND2X7 U17382 ( .A(n4280), .B(n4271), .Z(n3326) );
  HS65_LL_NAND2X7 U17383 ( .A(n9028), .B(n9046), .Z(n7676) );
  HS65_LL_NAND2X7 U17384 ( .A(n9086), .B(n9104), .Z(n7714) );
  HS65_LL_NAND2X7 U17385 ( .A(n1831), .B(n1842), .Z(n1555) );
  HS65_LL_NAND2X7 U17386 ( .A(n8986), .B(n8985), .Z(n8661) );
  HS65_LL_NAND2X7 U17387 ( .A(n5854), .B(n5855), .Z(n4923) );
  HS65_LL_NAND2X7 U17388 ( .A(n5913), .B(n5914), .Z(n4976) );
  HS65_LL_NAND2X7 U17389 ( .A(n7446), .B(n7447), .Z(n6516) );
  HS65_LL_NAND2X7 U17390 ( .A(n7505), .B(n7506), .Z(n6569) );
  HS65_LL_NAND2X7 U17391 ( .A(n8989), .B(n8967), .Z(n7861) );
  HS65_LL_NAND2X7 U17392 ( .A(n8986), .B(n8987), .Z(n7848) );
  HS65_LL_NAND2X7 U17393 ( .A(n5744), .B(n5745), .Z(n4566) );
  HS65_LL_NAND2X7 U17394 ( .A(n7336), .B(n7337), .Z(n6159) );
  HS65_LL_NAND2X7 U17395 ( .A(n8988), .B(n8968), .Z(n7992) );
  HS65_LL_NAND2X7 U17396 ( .A(n8907), .B(n8908), .Z(n8540) );
  HS65_LL_NAND2X7 U17397 ( .A(n4264), .B(n4281), .Z(n3141) );
  HS65_LL_NAND2X7 U17398 ( .A(n5740), .B(n5739), .Z(n4710) );
  HS65_LL_NAND2X7 U17399 ( .A(n7332), .B(n7331), .Z(n6303) );
  HS65_LL_NAND2X7 U17400 ( .A(n5802), .B(n5810), .Z(n4533) );
  HS65_LL_NAND2X7 U17401 ( .A(n7394), .B(n7402), .Z(n6126) );
  HS65_LL_NAND2X7 U17402 ( .A(n5863), .B(n5864), .Z(n4586) );
  HS65_LL_NAND2X7 U17403 ( .A(n7514), .B(n7515), .Z(n6196) );
  HS65_LL_NAND2X7 U17404 ( .A(n7457), .B(n7458), .Z(n6179) );
  HS65_LL_NAND2X7 U17405 ( .A(n5922), .B(n5923), .Z(n4603) );
  HS65_LL_NAND2X7 U17406 ( .A(n4266), .B(n4265), .Z(n3692) );
  HS65_LL_NAND2X7 U17407 ( .A(n9102), .B(n9077), .Z(n7874) );
  HS65_LL_NAND2X7 U17408 ( .A(n9044), .B(n9019), .Z(n7835) );
  HS65_LL_NAND2X7 U17409 ( .A(n9048), .B(n9027), .Z(n7619) );
  HS65_LL_NAND2X7 U17410 ( .A(n9106), .B(n9085), .Z(n7656) );
  HS65_LL_NAND2X7 U17411 ( .A(n8979), .B(n8990), .Z(n7750) );
  HS65_LL_NAND2X7 U17412 ( .A(n4211), .B(n4212), .Z(n3491) );
  HS65_LL_NAND2X7 U17413 ( .A(n2583), .B(n2604), .Z(n2274) );
  HS65_LL_NAND2X7 U17414 ( .A(n1455), .B(n1476), .Z(n1146) );
  HS65_LL_NAND2X7 U17415 ( .A(n2207), .B(n2228), .Z(n1898) );
  HS65_LL_NAND2X7 U17416 ( .A(n8931), .B(n8917), .Z(n8871) );
  HS65_LL_NAND2X7 U17417 ( .A(n4328), .B(n4329), .Z(n2832) );
  HS65_LL_NAND2X7 U17418 ( .A(n5874), .B(n5870), .Z(n4748) );
  HS65_LL_NAND2X7 U17419 ( .A(n5933), .B(n5929), .Z(n4774) );
  HS65_LL_NAND2X7 U17420 ( .A(n7461), .B(n7453), .Z(n6328) );
  HS65_LL_NAND2X7 U17421 ( .A(n7525), .B(n7521), .Z(n6367) );
  HS65_LL_NAND2X7 U17422 ( .A(n1831), .B(n1852), .Z(n1522) );
  HS65_LL_NAND2X7 U17423 ( .A(n5862), .B(n5852), .Z(n4747) );
  HS65_LL_NAND2X7 U17424 ( .A(n5921), .B(n5911), .Z(n4773) );
  HS65_LL_NAND2X7 U17425 ( .A(n7455), .B(n7444), .Z(n6327) );
  HS65_LL_NAND2X7 U17426 ( .A(n7513), .B(n7503), .Z(n6366) );
  HS65_LL_NAND2X7 U17427 ( .A(n5933), .B(n5911), .Z(n5554) );
  HS65_LL_NAND2X7 U17428 ( .A(n7525), .B(n7503), .Z(n7146) );
  HS65_LL_NAND2X7 U17429 ( .A(n5874), .B(n5852), .Z(n5532) );
  HS65_LL_NAND2X7 U17430 ( .A(n7461), .B(n7444), .Z(n7124) );
  HS65_LL_NAND2X7 U17431 ( .A(n7401), .B(n7382), .Z(n7171) );
  HS65_LL_NAND2X7 U17432 ( .A(n5809), .B(n5790), .Z(n5579) );
  HS65_LL_NAND2X7 U17433 ( .A(n8970), .B(n8971), .Z(n7981) );
  HS65_LL_NOR2X6 U17434 ( .A(n181), .B(n176), .Z(n4158) );
  HS65_LL_NOR2X6 U17435 ( .A(n486), .B(n487), .Z(n5930) );
  HS65_LL_NOR2X6 U17436 ( .A(n269), .B(n270), .Z(n5871) );
  HS65_LL_NOR2X6 U17437 ( .A(n311), .B(n312), .Z(n7522) );
  HS65_LL_NOR2X6 U17438 ( .A(n43), .B(n48), .Z(n5751) );
  HS65_LL_NOR2X6 U17439 ( .A(n698), .B(n703), .Z(n5813) );
  HS65_LL_NOR2X6 U17440 ( .A(n522), .B(n527), .Z(n7405) );
  HS65_LL_NOR2X6 U17441 ( .A(n565), .B(n570), .Z(n7343) );
  HS65_LL_NOR2X6 U17442 ( .A(n87), .B(n92), .Z(n7466) );
  HS65_LL_NAND2X7 U17443 ( .A(n5740), .B(n5748), .Z(n4477) );
  HS65_LL_NAND2X7 U17444 ( .A(n7332), .B(n7340), .Z(n6070) );
  HS65_LL_NAND2X7 U17445 ( .A(n4272), .B(n4282), .Z(n2970) );
  HS65_LLS_XOR2X6 U17446 ( .A(n2279), .B(n946), .Z(n1003) );
  HS65_LL_NOR3X4 U17447 ( .A(n2280), .B(n2281), .C(n2282), .Z(n2279) );
  HS65_LL_OAI212X5 U17448 ( .A(n2283), .B(n2284), .C(n2285), .D(n2238), .E(
        n2286), .Z(n2282) );
  HS65_LL_NAND4ABX3 U17449 ( .A(n2292), .B(n2293), .C(n2294), .D(n2295), .Z(
        n2281) );
  HS65_LLS_XOR2X6 U17450 ( .A(n1527), .B(n955), .Z(n987) );
  HS65_LL_NOR3X4 U17451 ( .A(n1528), .B(n1529), .C(n1530), .Z(n1527) );
  HS65_LL_OAI212X5 U17452 ( .A(n1531), .B(n1532), .C(n1533), .D(n1486), .E(
        n1534), .Z(n1530) );
  HS65_LL_NAND4ABX3 U17453 ( .A(n1540), .B(n1541), .C(n1542), .D(n1543), .Z(
        n1529) );
  HS65_LL_NAND2X7 U17454 ( .A(n4267), .B(n4270), .Z(n3731) );
  HS65_LL_NAND2X7 U17455 ( .A(n4331), .B(n4339), .Z(n2995) );
  HS65_LL_NAND2X7 U17456 ( .A(n4215), .B(n4210), .Z(n2857) );
  HS65_LLS_XOR2X6 U17457 ( .A(n2126), .B(n947), .Z(n998) );
  HS65_LL_NOR4ABX2 U17458 ( .A(n2127), .B(n2128), .C(n2129), .D(n2130), .Z(
        n2126) );
  HS65_LL_CBI4I1X5 U17459 ( .A(n1915), .B(n1863), .C(n1897), .D(n2093), .Z(
        n2130) );
  HS65_LL_AOI212X4 U17460 ( .A(n770), .B(n789), .C(n778), .D(n1875), .E(n2145), 
        .Z(n2128) );
  HS65_LLS_XOR2X6 U17461 ( .A(n1750), .B(n952), .Z(n990) );
  HS65_LL_NOR4ABX2 U17462 ( .A(n1751), .B(n1752), .C(n1753), .D(n1754), .Z(
        n1750) );
  HS65_LL_CBI4I1X5 U17463 ( .A(n1539), .B(n1487), .C(n1521), .D(n1717), .Z(
        n1754) );
  HS65_LL_AOI212X4 U17464 ( .A(n811), .B(n830), .C(n819), .D(n1499), .E(n1769), 
        .Z(n1752) );
  HS65_LLS_XOR2X6 U17465 ( .A(n1857), .B(n949), .Z(n993) );
  HS65_LL_NOR3X4 U17466 ( .A(n1858), .B(n1859), .C(n1860), .Z(n1857) );
  HS65_LL_NAND4ABX3 U17467 ( .A(n1871), .B(n1872), .C(n1873), .D(n1874), .Z(
        n1859) );
  HS65_LL_OAI212X5 U17468 ( .A(n1861), .B(n1862), .C(n1863), .D(n1864), .E(
        n1865), .Z(n1860) );
  HS65_LLS_XOR2X6 U17469 ( .A(n2321), .B(n945), .Z(n1004) );
  HS65_LL_NOR3X4 U17470 ( .A(n2322), .B(n2323), .C(n2324), .Z(n2321) );
  HS65_LL_OAI212X5 U17471 ( .A(n2325), .B(n2240), .C(n2326), .D(n2327), .E(
        n2328), .Z(n2324) );
  HS65_LL_NAND4ABX3 U17472 ( .A(n2329), .B(n2330), .C(n2331), .D(n2332), .Z(
        n2323) );
  HS65_LLS_XOR2X6 U17473 ( .A(n1569), .B(n954), .Z(n988) );
  HS65_LL_NOR3X4 U17474 ( .A(n1570), .B(n1571), .C(n1572), .Z(n1569) );
  HS65_LL_NAND4ABX3 U17475 ( .A(n1577), .B(n1578), .C(n1579), .D(n1580), .Z(
        n1571) );
  HS65_LL_OAI212X5 U17476 ( .A(n1573), .B(n1488), .C(n1574), .D(n1575), .E(
        n1576), .Z(n1572) );
  HS65_LLS_XOR2X6 U17477 ( .A(n948), .B(n1884), .Z(n994) );
  HS65_LL_NAND4ABX3 U17478 ( .A(n1885), .B(n1886), .C(n1887), .D(n1888), .Z(
        n1884) );
  HS65_LL_AOI212X4 U17479 ( .A(n791), .B(n757), .C(n788), .D(n769), .E(n1894), 
        .Z(n1887) );
  HS65_LL_CBI4I1X5 U17480 ( .A(n1896), .B(n1897), .C(n1898), .D(n1899), .Z(
        n1886) );
  HS65_LLS_XOR2X6 U17481 ( .A(n943), .B(n2524), .Z(n1007) );
  HS65_LL_NAND4ABX3 U17482 ( .A(n2525), .B(n2526), .C(n2527), .D(n2528), .Z(
        n2524) );
  HS65_LL_CB4I6X9 U17483 ( .A(n885), .B(n890), .C(n912), .D(n2462), .Z(n2525)
         );
  HS65_LL_AOI222X2 U17484 ( .A(n904), .B(n882), .C(n901), .D(n2547), .E(n913), 
        .F(n881), .Z(n2527) );
  HS65_LLS_XOR2X6 U17485 ( .A(n951), .B(n1772), .Z(n991) );
  HS65_LL_NAND4ABX3 U17486 ( .A(n1773), .B(n1774), .C(n1775), .D(n1776), .Z(
        n1772) );
  HS65_LL_AOI222X2 U17487 ( .A(n822), .B(n800), .C(n819), .D(n1795), .E(n831), 
        .F(n799), .Z(n1775) );
  HS65_LL_CB4I6X9 U17488 ( .A(n803), .B(n808), .C(n830), .D(n1710), .Z(n1773)
         );
  HS65_LLS_XOR2X6 U17489 ( .A(n950), .B(n1797), .Z(n992) );
  HS65_LL_NAND4ABX3 U17490 ( .A(n1798), .B(n1799), .C(n1800), .D(n1801), .Z(
        n1797) );
  HS65_LL_MX41X7 U17491 ( .D0(n811), .S0(n828), .D1(n812), .S1(n820), .D2(n831), .S2(n804), .D3(n832), .S3(n1561), .Z(n1799) );
  HS65_LL_NOR4ABX2 U17492 ( .A(n1559), .B(n1694), .C(n1802), .D(n1708), .Z(
        n1801) );
  HS65_LL_NAND2X7 U17493 ( .A(n5910), .B(n5911), .Z(n4995) );
  HS65_LL_NAND2X7 U17494 ( .A(n7502), .B(n7503), .Z(n6588) );
  HS65_LL_NAND2X7 U17495 ( .A(n7443), .B(n7444), .Z(n6476) );
  HS65_LL_NAND2X7 U17496 ( .A(n5855), .B(n5876), .Z(n4882) );
  HS65_LL_NAND2X7 U17497 ( .A(n5914), .B(n5935), .Z(n4994) );
  HS65_LL_NAND2X7 U17498 ( .A(n7506), .B(n7527), .Z(n6587) );
  HS65_LL_NAND2X7 U17499 ( .A(n7447), .B(n7469), .Z(n6475) );
  HS65_LLS_XOR2X6 U17500 ( .A(n938), .B(n983), .Z(n1079) );
  HS65_LLS_XOR2X6 U17501 ( .A(n941), .B(n978), .Z(n1074) );
  HS65_LL_NAND2X7 U17502 ( .A(n5924), .B(n5923), .Z(n5382) );
  HS65_LL_NAND2X7 U17503 ( .A(n5865), .B(n5864), .Z(n5267) );
  HS65_LL_NAND2X7 U17504 ( .A(n7516), .B(n7515), .Z(n6974) );
  HS65_LL_NAND2X7 U17505 ( .A(n7459), .B(n7458), .Z(n6859) );
  HS65_LL_NAND2X7 U17506 ( .A(n5744), .B(n5739), .Z(n4478) );
  HS65_LL_NAND2X7 U17507 ( .A(n7336), .B(n7331), .Z(n6071) );
  HS65_LL_NAND2X7 U17508 ( .A(n7398), .B(n7393), .Z(n6127) );
  HS65_LL_NAND2X7 U17509 ( .A(n5865), .B(n5855), .Z(n4454) );
  HS65_LL_NAND2X7 U17510 ( .A(n7516), .B(n7506), .Z(n6086) );
  HS65_LL_NAND2X7 U17511 ( .A(n7459), .B(n7447), .Z(n6047) );
  HS65_LL_NAND2X7 U17512 ( .A(n5924), .B(n5914), .Z(n4493) );
  HS65_LLS_XOR2X6 U17513 ( .A(n944), .B(n2383), .Z(n1005) );
  HS65_LL_NAND4ABX3 U17514 ( .A(n2384), .B(n2385), .C(n2386), .D(n2387), .Z(
        n2383) );
  HS65_LL_MX41X7 U17515 ( .D0(n906), .S0(n884), .D1(n908), .S1(n891), .D2(n901), .S2(n894), .D3(n885), .S3(n915), .Z(n2384) );
  HS65_LL_AOI212X4 U17516 ( .A(n896), .B(n2388), .C(n912), .D(n2365), .E(n2389), .Z(n2387) );
  HS65_LLS_XOR2X6 U17517 ( .A(n953), .B(n1631), .Z(n989) );
  HS65_LL_NAND4ABX3 U17518 ( .A(n1632), .B(n1633), .C(n1634), .D(n1635), .Z(
        n1631) );
  HS65_LL_MX41X7 U17519 ( .D0(n801), .S0(n825), .D1(n829), .S1(n813), .D2(n799), .S2(n820), .D3(n831), .S3(n1561), .Z(n1633) );
  HS65_LL_AOI212X4 U17520 ( .A(n814), .B(n1636), .C(n830), .D(n1613), .E(n1637), .Z(n1635) );
  HS65_LLS_XOR3X2 U17521 ( .A(n2759), .B(n938), .C(n2806), .Z(n5966) );
  HS65_LLS_XOR3X2 U17522 ( .A(n2767), .B(n957), .C(n2814), .Z(n4373) );
  HS65_LL_NAND2X7 U17523 ( .A(n4151), .B(n4140), .Z(n2917) );
  HS65_LL_NAND2X7 U17524 ( .A(n5805), .B(n5789), .Z(n5148) );
  HS65_LL_NAND2X7 U17525 ( .A(n4147), .B(n4148), .Z(n3033) );
  HS65_LL_NAND2X7 U17526 ( .A(n5812), .B(n5813), .Z(n5572) );
  HS65_LL_NAND2X7 U17527 ( .A(n5810), .B(n5814), .Z(n5135) );
  HS65_LL_NAND2X7 U17528 ( .A(n7402), .B(n7406), .Z(n6727) );
  HS65_LL_NAND2X7 U17529 ( .A(n4153), .B(n4155), .Z(n3043) );
  HS65_LL_NAND2X7 U17530 ( .A(n4157), .B(n4158), .Z(n3574) );
  HS65_LL_NAND2X7 U17531 ( .A(n4150), .B(n4152), .Z(n3032) );
  HS65_LL_NAND2X7 U17532 ( .A(n4140), .B(n4154), .Z(n3270) );
  HS65_LL_NAND2X7 U17533 ( .A(n4145), .B(n4157), .Z(n4093) );
  HS65_LL_NAND2X7 U17534 ( .A(n9045), .B(n9040), .Z(n8005) );
  HS65_LL_NAND2X7 U17535 ( .A(n4159), .B(n4150), .Z(n3225) );
  HS65_LL_NAND2X7 U17536 ( .A(n4137), .B(n4138), .Z(n3252) );
  HS65_LL_NAND2X7 U17537 ( .A(n4138), .B(n4150), .Z(n3053) );
  HS65_LL_NAND2X7 U17538 ( .A(n4147), .B(n4153), .Z(n3982) );
  HS65_LL_NAND2X7 U17539 ( .A(n4137), .B(n4140), .Z(n2914) );
  HS65_LL_NAND2X7 U17540 ( .A(n9103), .B(n9100), .Z(n7870) );
  HS65_LL_NAND2X7 U17541 ( .A(n5812), .B(n5789), .Z(n4848) );
  HS65_LL_NAND2X7 U17542 ( .A(n7404), .B(n7381), .Z(n6441) );
  HS65_LL_NAND2X7 U17543 ( .A(n4159), .B(n4137), .Z(n3286) );
  HS65_LL_NAND2X7 U17544 ( .A(n9047), .B(n9049), .Z(n7632) );
  HS65_LL_NAND2X7 U17545 ( .A(n9105), .B(n9107), .Z(n7652) );
  HS65_LL_IVX9 U17546 ( .A(n968), .Z(n963) );
  HS65_LL_NAND2X7 U17547 ( .A(n4157), .B(n4148), .Z(n3251) );
  HS65_LL_NAND2X7 U17548 ( .A(n5750), .B(n5727), .Z(n4709) );
  HS65_LL_NAND2X7 U17549 ( .A(n7342), .B(n7319), .Z(n6302) );
  HS65_LL_NAND2X7 U17550 ( .A(n4146), .B(n4153), .Z(n3034) );
  HS65_LL_NAND2X7 U17551 ( .A(n7395), .B(n7392), .Z(n6118) );
  HS65_LL_NAND2X7 U17552 ( .A(n5803), .B(n5800), .Z(n4525) );
  HS65_LL_NAND2X7 U17553 ( .A(n5743), .B(n5727), .Z(n5026) );
  HS65_LL_NAND2X7 U17554 ( .A(n7335), .B(n7319), .Z(n6619) );
  HS65_LL_NAND2X7 U17555 ( .A(n5803), .B(n5814), .Z(n4809) );
  HS65_LL_NAND2X7 U17556 ( .A(n7395), .B(n7406), .Z(n6402) );
  HS65_LL_NAND2X7 U17557 ( .A(n5802), .B(n5801), .Z(n4847) );
  HS65_LL_NAND2X7 U17558 ( .A(n7394), .B(n7393), .Z(n6440) );
  HS65_LL_NAND2X7 U17559 ( .A(n4203), .B(n4220), .Z(n3114) );
  HS65_LL_NAND2X7 U17560 ( .A(n971), .B(n966), .Z(n972) );
  HS65_LL_NAND2X7 U17561 ( .A(n9019), .B(n9034), .Z(n7620) );
  HS65_LL_NAND2X7 U17562 ( .A(n9077), .B(n9092), .Z(n7660) );
  HS65_LL_NAND2X7 U17563 ( .A(n4151), .B(n4152), .Z(n3615) );
  HS65_LL_NAND2X7 U17564 ( .A(n5800), .B(n5801), .Z(n4849) );
  HS65_LL_NAND2X7 U17565 ( .A(n7392), .B(n7393), .Z(n6442) );
  HS65_LL_NAND2X7 U17566 ( .A(n5747), .B(n5743), .Z(n4551) );
  HS65_LL_NAND2X7 U17567 ( .A(n7339), .B(n7335), .Z(n6144) );
  HS65_LL_NAND2X7 U17568 ( .A(n4146), .B(n4148), .Z(n3269) );
  HS65_LL_NAND2X7 U17569 ( .A(n9100), .B(n9086), .Z(n7920) );
  HS65_LL_NAND2X7 U17570 ( .A(n9042), .B(n9028), .Z(n7822) );
  HS65_LL_NAND2X7 U17571 ( .A(\u0/r0/N80 ), .B(n966), .Z(n967) );
  HS65_LL_NAND2X7 U17572 ( .A(n4159), .B(n4154), .Z(n3271) );
  HS65_LL_NAND2X7 U17573 ( .A(n5745), .B(n5752), .Z(n5472) );
  HS65_LL_NAND2X7 U17574 ( .A(n7337), .B(n7344), .Z(n7064) );
  HS65_LL_NAND2X7 U17575 ( .A(n4138), .B(n4154), .Z(n3047) );
  HS65_LL_NAND2X7 U17576 ( .A(n5809), .B(n5805), .Z(n4628) );
  HS65_LL_NAND2X7 U17577 ( .A(n7401), .B(n7397), .Z(n6221) );
  HS65_LL_NAND2X7 U17578 ( .A(n4145), .B(n4147), .Z(n2915) );
  HS65_LL_NAND2X7 U17579 ( .A(n5789), .B(n5790), .Z(n4627) );
  HS65_LL_NAND2X7 U17580 ( .A(n7381), .B(n7382), .Z(n6220) );
  HS65_LL_NAND2X7 U17581 ( .A(n9100), .B(n9106), .Z(n8168) );
  HS65_LL_NAND2X7 U17582 ( .A(n9042), .B(n9048), .Z(n8145) );
  HS65_LL_NAND2X7 U17583 ( .A(n4145), .B(n4155), .Z(n3984) );
  HS65_LL_NAND2X7 U17584 ( .A(n5738), .B(n5739), .Z(n4711) );
  HS65_LL_NAND2X7 U17585 ( .A(n7330), .B(n7331), .Z(n6304) );
  HS65_LL_IVX9 U17586 ( .A(n2610), .Z(n1) );
  HS65_LL_OAI311X5 U17587 ( .A(n972), .B(n964), .C(n963), .D(n973), .E(n9145), 
        .Z(\u0/r0/N70 ) );
  HS65_LL_NAND3X5 U17588 ( .A(n9145), .B(n964), .C(n974), .Z(n969) );
  HS65_LL_NAND2X7 U17589 ( .A(n5851), .B(n5852), .Z(n4883) );
  HS65_LL_NAND2X7 U17590 ( .A(n7396), .B(n7382), .Z(n6462) );
  HS65_LL_NAND2X7 U17591 ( .A(n5804), .B(n5790), .Z(n4869) );
  HS65_LL_NOR3AX2 U17592 ( .A(n971), .B(n963), .C(n966), .Z(n974) );
  HS65_LL_NAND2X7 U17593 ( .A(n7393), .B(n7406), .Z(n6461) );
  HS65_LL_NAND2X7 U17594 ( .A(n5801), .B(n5814), .Z(n4868) );
  HS65_LL_NAND2X7 U17595 ( .A(n5739), .B(n5752), .Z(n4667) );
  HS65_LL_NAND2X7 U17596 ( .A(n7331), .B(n7344), .Z(n6260) );
  HS65_LL_NAND2X7 U17597 ( .A(n5806), .B(n5810), .Z(n5150) );
  HS65_LL_NAND2X7 U17598 ( .A(n7398), .B(n7402), .Z(n6742) );
  HS65_LL_NAND2X7 U17599 ( .A(n5806), .B(n5801), .Z(n4534) );
  HS65_LL_NAND2X7 U17600 ( .A(n5744), .B(n5748), .Z(n5028) );
  HS65_LL_NAND2X7 U17601 ( .A(n7336), .B(n7340), .Z(n6621) );
  HS65_LL_OAI31X5 U17602 ( .A(n963), .B(n964), .C(n967), .D(n970), .Z(
        \u0/r0/N74 ) );
  HS65_LL_OAI31X5 U17603 ( .A(n706), .B(n964), .C(n972), .D(n969), .Z(
        \u0/r0/N72 ) );
  HS65_LL_NOR2X6 U17604 ( .A(n5), .B(n1), .Z(n2611) );
  HS65_LL_OAI31X5 U17605 ( .A(n707), .B(n972), .C(n963), .D(n970), .Z(
        \u0/r0/N71 ) );
  HS65_LL_IVX9 U17606 ( .A(\u0/r0/N78 ), .Z(n707) );
  HS65_LL_NOR3X4 U17607 ( .A(n967), .B(n968), .C(n964), .Z(\u0/r0/N76 ) );
  HS65_LLS_XNOR2X6 U17608 ( .A(n2708), .B(n817), .Z(N471) );
  HS65_LLS_XNOR2X6 U17609 ( .A(n2631), .B(n919), .Z(N403) );
  HS65_LLS_XNOR2X6 U17610 ( .A(n2687), .B(n837), .Z(N467) );
  HS65_LLS_XNOR2X6 U17611 ( .A(n2638), .B(n918), .Z(N404) );
  HS65_LLS_XNOR2X6 U17612 ( .A(n2692), .B(n836), .Z(N468) );
  HS65_LLS_XNOR2X6 U17613 ( .A(n2713), .B(n816), .Z(N472) );
  HS65_LLS_XNOR2X6 U17614 ( .A(n2703), .B(n818), .Z(N470) );
  HS65_LL_NOR2X6 U17615 ( .A(n968), .B(n9138), .Z(\u0/r0/N79 ) );
  HS65_LL_NOR2X6 U17616 ( .A(n971), .B(n9137), .Z(\u0/r0/N80 ) );
  HS65_LLS_XNOR2X6 U17617 ( .A(n2682), .B(n920), .Z(N402) );
  HS65_LLS_XNOR2X6 U17618 ( .A(n2698), .B(n835), .Z(N469) );
  HS65_LLS_XNOR2X6 U17619 ( .A(n2645), .B(n917), .Z(N405) );
  HS65_LLS_XNOR2X6 U17620 ( .A(n2672), .B(n856), .Z(N441) );
  HS65_LLS_XNOR2X6 U17621 ( .A(n2674), .B(n897), .Z(N409) );
  HS65_LLS_XNOR2X6 U17622 ( .A(n2718), .B(n815), .Z(N473) );
  HS65_LLS_XNOR2X6 U17623 ( .A(n2673), .B(n775), .Z(N504) );
  HS65_LLS_XNOR2X6 U17624 ( .A(n2652), .B(n900), .Z(N406) );
  HS65_LLS_XNOR2X6 U17625 ( .A(n2630), .B(n879), .Z(N434) );
  HS65_LLS_XNOR2X6 U17626 ( .A(n2722), .B(n797), .Z(N498) );
  HS65_LLS_XNOR2X6 U17627 ( .A(n3533), .B(n962), .Z(N378) );
  HS65_LLS_XNOR2X6 U17628 ( .A(n3208), .B(n942), .Z(N386) );
  HS65_LLS_XNOR2X6 U17629 ( .A(n2769), .B(n944), .Z(N478) );
  HS65_LLS_XNOR2X6 U17630 ( .A(n2771), .B(n946), .Z(N476) );
  HS65_LLS_XNOR2X6 U17631 ( .A(n3002), .B(n930), .Z(N397) );
  HS65_LLS_XNOR2X6 U17632 ( .A(n2819), .B(n955), .Z(N412) );
  HS65_LLS_XNOR2X6 U17633 ( .A(n3212), .B(n959), .Z(N382) );
  HS65_LLS_XNOR2X6 U17634 ( .A(n3007), .B(n938), .Z(N392) );
  HS65_LLS_XNOR2X6 U17635 ( .A(n3210), .B(n957), .Z(N384) );
  HS65_LLS_XNOR2X6 U17636 ( .A(n3000), .B(n928), .Z(N399) );
  HS65_LLS_XNOR2X6 U17637 ( .A(n2816), .B(n952), .Z(N415) );
  HS65_LLS_XNOR2X6 U17638 ( .A(n2815), .B(n951), .Z(N416) );
  HS65_LLS_XNOR2X6 U17639 ( .A(n3209), .B(n956), .Z(N385) );
  HS65_LLS_XNOR2X6 U17640 ( .A(n2814), .B(n950), .Z(N417) );
  HS65_LLS_XNOR2X6 U17641 ( .A(n3207), .B(n941), .Z(N387) );
  HS65_LLS_XNOR2X6 U17642 ( .A(n2792), .B(n947), .Z(N447) );
  HS65_LLS_XNOR2X6 U17643 ( .A(n2784), .B(n933), .Z(N455) );
  HS65_LLS_XNOR2X6 U17644 ( .A(n2789), .B(n934), .Z(N450) );
  HS65_LLS_XNOR2X6 U17645 ( .A(n2797), .B(n949), .Z(N442) );
  HS65_LLS_XNOR2X6 U17646 ( .A(n3213), .B(n960), .Z(N381) );
  HS65_LLS_XNOR2X6 U17647 ( .A(n2817), .B(n953), .Z(N414) );
  HS65_LLS_XNOR2X6 U17648 ( .A(n2818), .B(n954), .Z(N413) );
  HS65_LLS_XNOR2X6 U17649 ( .A(n3004), .B(n931), .Z(N395) );
  HS65_LLS_XNOR2X6 U17650 ( .A(n3532), .B(n961), .Z(N379) );
  HS65_LLS_XNOR2X6 U17651 ( .A(n3008), .B(n939), .Z(N391) );
  HS65_LLS_XNOR2X6 U17652 ( .A(n3211), .B(n958), .Z(N383) );
  HS65_LL_IVX9 U17653 ( .A(n2613), .Z(n705) );
  HS65_LL_OA12X9 U17654 ( .A(n9142), .B(n973), .C(n969), .Z(n970) );
  HS65_LL_BFX9 U17655 ( .A(n9136), .Z(n9135) );
  HS65_LL_NOR2X6 U17656 ( .A(n9138), .B(n966), .Z(\u0/r0/N81 ) );
  HS65_LL_IVX9 U17657 ( .A(n9150), .Z(n9149) );
  HS65_LLS_XNOR3X2 U17658 ( .A(n1151), .B(\u0/rcon [29]), .C(w0[29]), .Z(n979)
         );
  HS65_LL_NOR3X4 U17659 ( .A(n1152), .B(n1153), .C(n1154), .Z(n1151) );
  HS65_LL_OAI212X5 U17660 ( .A(n1155), .B(n1156), .C(n1157), .D(n1110), .E(
        n1158), .Z(n1154) );
  HS65_LL_NAND4ABX3 U17661 ( .A(n1164), .B(n1165), .C(n1166), .D(n1167), .Z(
        n1153) );
  HS65_LL_NOR2X6 U17662 ( .A(w3[3]), .B(w3[2]), .Z(n2229) );
  HS65_LL_NOR2X6 U17663 ( .A(w3[19]), .B(w3[18]), .Z(n1477) );
  HS65_LL_NOR2X6 U17664 ( .A(n775), .B(w3[0]), .Z(n2209) );
  HS65_LL_NOR2X6 U17665 ( .A(n337), .B(sa02[4]), .Z(n8928) );
  HS65_LL_NOR2X6 U17666 ( .A(n381), .B(sa31[4]), .Z(n8977) );
  HS65_LL_NOR2X6 U17667 ( .A(sa31[7]), .B(sa31[6]), .Z(n8967) );
  HS65_LL_NOR2X6 U17668 ( .A(sa02[7]), .B(sa02[6]), .Z(n8907) );
  HS65_LL_NOR2X6 U17669 ( .A(w3[27]), .B(w3[26]), .Z(n2605) );
  HS65_LL_NOR2X6 U17670 ( .A(n836), .B(w3[12]), .Z(n1855) );
  HS65_LL_NOR2X6 U17671 ( .A(n918), .B(w3[28]), .Z(n2607) );
  HS65_LL_NOR2X6 U17672 ( .A(n898), .B(w3[24]), .Z(n2585) );
  HS65_LL_NOR2X6 U17673 ( .A(n857), .B(w3[16]), .Z(n1457) );
  HS65_LL_NOR2X6 U17674 ( .A(n816), .B(w3[8]), .Z(n1833) );
  HS65_LL_NOR2X6 U17675 ( .A(n877), .B(w3[20]), .Z(n1479) );
  HS65_LL_NOR2X6 U17676 ( .A(n795), .B(w3[4]), .Z(n2231) );
  HS65_LL_NOR2X6 U17677 ( .A(w3[11]), .B(w3[10]), .Z(n1853) );
  HS65_LL_NOR2X6 U17678 ( .A(sa21[3]), .B(sa21[2]), .Z(n4340) );
  HS65_LL_NOR2X6 U17679 ( .A(sa32[3]), .B(sa32[2]), .Z(n4221) );
  HS65_LL_NOR2X6 U17680 ( .A(sa02[3]), .B(sa02[2]), .Z(n8910) );
  HS65_LL_NOR2X6 U17681 ( .A(sa31[3]), .B(sa31[2]), .Z(n8970) );
  HS65_LL_NOR2X6 U17682 ( .A(n401), .B(sa31[2]), .Z(n8992) );
  HS65_LL_NOR2X6 U17683 ( .A(n357), .B(sa02[2]), .Z(n8924) );
  HS65_LL_NOR2X6 U17684 ( .A(n859), .B(w3[18]), .Z(n1466) );
  HS65_LL_NOR2X6 U17685 ( .A(n777), .B(w3[2]), .Z(n2218) );
  HS65_LL_NOR2X6 U17686 ( .A(n837), .B(w3[15]), .Z(n1854) );
  HS65_LL_NOR2X6 U17687 ( .A(n876), .B(w3[21]), .Z(n1474) );
  HS65_LL_NOR2X6 U17688 ( .A(n794), .B(w3[5]), .Z(n2226) );
  HS65_LL_NOR2X6 U17689 ( .A(n43), .B(sa33[2]), .Z(n5727) );
  HS65_LL_NOR2X6 U17690 ( .A(n565), .B(sa30[2]), .Z(n7319) );
  HS65_LL_NOR2X6 U17691 ( .A(n116), .B(sa13[4]), .Z(n9102) );
  HS65_LL_NOR2X6 U17692 ( .A(n596), .B(sa20[4]), .Z(n9044) );
  HS65_LL_NOR2X6 U17693 ( .A(n133), .B(sa13[2]), .Z(n9100) );
  HS65_LL_NOR2X6 U17694 ( .A(n613), .B(sa20[2]), .Z(n9042) );
  HS65_LL_NOR2X6 U17695 ( .A(sa21[7]), .B(sa21[6]), .Z(n4328) );
  HS65_LL_NOR2X6 U17696 ( .A(n161), .B(sa03[4]), .Z(n4159) );
  HS65_LL_NOR2X6 U17697 ( .A(n597), .B(sa20[5]), .Z(n9047) );
  HS65_LL_NOR2X6 U17698 ( .A(n117), .B(sa13[5]), .Z(n9105) );
  HS65_LL_NOR2X6 U17699 ( .A(n114), .B(sa13[6]), .Z(n9109) );
  HS65_LL_NOR2X6 U17700 ( .A(n594), .B(sa20[6]), .Z(n9051) );
  HS65_LL_NOR2X6 U17701 ( .A(n206), .B(sa32[4]), .Z(n4218) );
  HS65_LL_NOR2X6 U17702 ( .A(n269), .B(sa22[2]), .Z(n5862) );
  HS65_LL_NOR2X6 U17703 ( .A(n486), .B(sa11[2]), .Z(n5921) );
  HS65_LL_NOR2X6 U17704 ( .A(n698), .B(sa00[2]), .Z(n5789) );
  HS65_LL_NOR2X6 U17705 ( .A(n424), .B(sa21[4]), .Z(n4342) );
  HS65_LL_NOR2X6 U17706 ( .A(n642), .B(sa10[4]), .Z(n4278) );
  HS65_LL_NOR2X6 U17707 ( .A(sa02[1]), .B(sa02[0]), .Z(n8911) );
  HS65_LL_NOR2X6 U17708 ( .A(n87), .B(sa23[2]), .Z(n7455) );
  HS65_LL_NOR2X6 U17709 ( .A(n311), .B(sa12[2]), .Z(n7513) );
  HS65_LL_NOR2X6 U17710 ( .A(n522), .B(sa01[2]), .Z(n7381) );
  HS65_LL_NOR2X6 U17711 ( .A(n445), .B(sa21[0]), .Z(n4324) );
  HS65_LL_NOR2X6 U17712 ( .A(n662), .B(sa10[2]), .Z(n4264) );
  HS65_LL_NOR2X6 U17713 ( .A(sa21[5]), .B(sa21[4]), .Z(n4327) );
  HS65_LL_NOR2X6 U17714 ( .A(sa32[5]), .B(sa32[4]), .Z(n4203) );
  HS65_LL_NOR2X6 U17715 ( .A(sa31[5]), .B(sa31[4]), .Z(n8979) );
  HS65_LL_NOR2X6 U17716 ( .A(sa02[5]), .B(sa02[4]), .Z(n8926) );
  HS65_LL_NOR2X6 U17717 ( .A(sa10[5]), .B(sa10[4]), .Z(n4268) );
  HS65_LL_NOR2X6 U17718 ( .A(n205), .B(sa32[7]), .Z(n4220) );
  HS65_LL_NOR2X6 U17719 ( .A(n423), .B(sa21[7]), .Z(n4341) );
  HS65_LL_NOR2X6 U17720 ( .A(n425), .B(sa21[5]), .Z(n4337) );
  HS65_LL_NOR2X6 U17721 ( .A(n162), .B(sa03[5]), .Z(n4138) );
  HS65_LL_NOR2X6 U17722 ( .A(n900), .B(w3[26]), .Z(n2594) );
  HS65_LL_NOR2X6 U17723 ( .A(n919), .B(w3[31]), .Z(n2606) );
  HS65_LL_NOR2X6 U17724 ( .A(n878), .B(w3[23]), .Z(n1478) );
  HS65_LL_NOR2X6 U17725 ( .A(n796), .B(w3[7]), .Z(n2230) );
  HS65_LL_NOR2X6 U17726 ( .A(n818), .B(w3[10]), .Z(n1842) );
  HS65_LL_NOR2X6 U17727 ( .A(n835), .B(w3[13]), .Z(n1850) );
  HS65_LL_NOR2X6 U17728 ( .A(n917), .B(w3[29]), .Z(n2602) );
  HS65_LL_NOR2X6 U17729 ( .A(n26), .B(sa33[7]), .Z(n5745) );
  HS65_LL_NOR2X6 U17730 ( .A(n548), .B(sa30[7]), .Z(n7337) );
  HS65_LL_NOR2X6 U17731 ( .A(n664), .B(sa10[0]), .Z(n4265) );
  HS65_LL_NOR2X6 U17732 ( .A(n222), .B(sa32[2]), .Z(n4213) );
  HS65_LL_NOR2X6 U17733 ( .A(n444), .B(sa21[2]), .Z(n4323) );
  HS65_LL_NOR2X6 U17734 ( .A(sa03[1]), .B(sa03[0]), .Z(n4146) );
  HS65_LL_NOR2X6 U17735 ( .A(n879), .B(w3[22]), .Z(n1464) );
  HS65_LL_NOR2X6 U17736 ( .A(n797), .B(w3[6]), .Z(n2216) );
  HS65_LL_NOR2X6 U17737 ( .A(w3[23]), .B(w3[22]), .Z(n1458) );
  HS65_LL_NOR2X6 U17738 ( .A(w3[7]), .B(w3[6]), .Z(n2210) );
  HS65_LL_NOR2X6 U17739 ( .A(n249), .B(sa22[5]), .Z(n5854) );
  HS65_LL_NOR2X6 U17740 ( .A(n466), .B(sa11[5]), .Z(n5913) );
  HS65_LL_NOR2X6 U17741 ( .A(n682), .B(sa00[5]), .Z(n5800) );
  HS65_LL_NOR2X6 U17742 ( .A(n71), .B(sa23[5]), .Z(n7446) );
  HS65_LL_NOR2X6 U17743 ( .A(n291), .B(sa12[5]), .Z(n7505) );
  HS65_LL_NOR2X6 U17744 ( .A(n506), .B(sa01[5]), .Z(n7392) );
  HS65_LL_NOR2X6 U17745 ( .A(w3[1]), .B(w3[0]), .Z(n2232) );
  HS65_LL_NOR2X6 U17746 ( .A(sa10[7]), .B(sa10[6]), .Z(n4269) );
  HS65_LL_NOR2X6 U17747 ( .A(n379), .B(sa31[6]), .Z(n8978) );
  HS65_LL_NOR2X6 U17748 ( .A(n204), .B(sa32[6]), .Z(n4211) );
  HS65_LL_NOR2X6 U17749 ( .A(n414), .B(sa21[6]), .Z(n4326) );
  HS65_LL_NOR2X6 U17750 ( .A(n632), .B(sa10[6]), .Z(n4267) );
  HS65_LL_NOR2X6 U17751 ( .A(n331), .B(sa02[6]), .Z(n8929) );
  HS65_LL_NOR2X6 U17752 ( .A(n181), .B(sa03[3]), .Z(n4145) );
  HS65_LL_NOR2X6 U17753 ( .A(sa13[7]), .B(sa13[6]), .Z(n9107) );
  HS65_LL_NOR2X6 U17754 ( .A(sa20[7]), .B(sa20[6]), .Z(n9049) );
  HS65_LL_NOR2X6 U17755 ( .A(sa03[7]), .B(sa03[6]), .Z(n4150) );
  HS65_LL_NOR2X6 U17756 ( .A(sa10[3]), .B(sa10[2]), .Z(n4283) );
  HS65_LL_NOR2X6 U17757 ( .A(n176), .B(sa03[2]), .Z(n4148) );
  HS65_LL_NOR2X6 U17758 ( .A(sa03[3]), .B(sa03[2]), .Z(n4153) );
  HS65_LL_NOR2X6 U17759 ( .A(n160), .B(sa03[7]), .Z(n4154) );
  HS65_LL_NOR2X6 U17760 ( .A(n336), .B(sa02[7]), .Z(n8919) );
  HS65_LL_NOR2X6 U17761 ( .A(n115), .B(sa13[7]), .Z(n9077) );
  HS65_LL_NOR2X6 U17762 ( .A(n595), .B(sa20[7]), .Z(n9019) );
  HS65_LL_NOR2X6 U17763 ( .A(n643), .B(sa10[5]), .Z(n4280) );
  HS65_LL_NOR2X6 U17764 ( .A(n380), .B(sa31[7]), .Z(n8990) );
  HS65_LL_NOR2X6 U17765 ( .A(n227), .B(sa32[0]), .Z(n4219) );
  HS65_LL_NOR2X6 U17766 ( .A(sa33[3]), .B(sa33[2]), .Z(n5747) );
  HS65_LL_NOR2X6 U17767 ( .A(sa30[3]), .B(sa30[2]), .Z(n7339) );
  HS65_LL_NOR2X6 U17768 ( .A(sa22[3]), .B(sa22[2]), .Z(n5874) );
  HS65_LL_NOR2X6 U17769 ( .A(sa11[3]), .B(sa11[2]), .Z(n5933) );
  HS65_LL_NOR2X6 U17770 ( .A(sa12[3]), .B(sa12[2]), .Z(n7525) );
  HS65_LL_NOR2X6 U17771 ( .A(sa01[3]), .B(sa01[2]), .Z(n7401) );
  HS65_LL_NOR2X6 U17772 ( .A(sa23[3]), .B(sa23[2]), .Z(n7461) );
  HS65_LL_NOR2X6 U17773 ( .A(n402), .B(sa31[0]), .Z(n8985) );
  HS65_LL_NOR2X6 U17774 ( .A(n382), .B(sa31[5]), .Z(n8968) );
  HS65_LL_NOR2X6 U17775 ( .A(n359), .B(sa02[1]), .Z(n8930) );
  HS65_LL_NOR2X6 U17776 ( .A(n403), .B(sa31[1]), .Z(n8991) );
  HS65_LL_NOR2X6 U17777 ( .A(n641), .B(sa10[7]), .Z(n4277) );
  HS65_LL_NOR2X6 U17778 ( .A(n207), .B(sa32[5]), .Z(n4201) );
  HS65_LL_OAI22X6 U17779 ( .A(n6011), .B(n9129), .C(n9123), .D(n6012), .Z(N183) );
  HS65_LLS_XNOR2X6 U17780 ( .A(w1[13]), .B(text_in_r[77]), .Z(n6011) );
  HS65_LLS_XNOR3X2 U17781 ( .A(n2811), .B(n6013), .C(n5982), .Z(n6012) );
  HS65_LLS_XOR3X2 U17782 ( .A(n2762), .B(w1[13]), .C(n2786), .Z(n6013) );
  HS65_LL_OAI22X6 U17783 ( .A(n4418), .B(n9133), .C(n9126), .D(n4419), .Z(N247) );
  HS65_LLS_XNOR2X6 U17784 ( .A(w0[13]), .B(text_in_r[109]), .Z(n4418) );
  HS65_LLS_XNOR3X2 U17785 ( .A(n2819), .B(n4420), .C(n4389), .Z(n4419) );
  HS65_LLS_XOR3X2 U17786 ( .A(n2770), .B(w0[13]), .C(n2794), .Z(n4420) );
  HS65_LL_NOR2X6 U17787 ( .A(sa20[5]), .B(sa20[4]), .Z(n9034) );
  HS65_LL_NOR2X6 U17788 ( .A(sa13[5]), .B(sa13[4]), .Z(n9092) );
  HS65_LL_NOR2X6 U17789 ( .A(sa33[1]), .B(sa33[0]), .Z(n5743) );
  HS65_LL_NOR2X6 U17790 ( .A(sa30[1]), .B(sa30[0]), .Z(n7335) );
  HS65_LL_NOR2X6 U17791 ( .A(sa11[7]), .B(sa11[6]), .Z(n5936) );
  HS65_LL_NOR2X6 U17792 ( .A(sa12[7]), .B(sa12[6]), .Z(n7528) );
  HS65_LL_NOR2X6 U17793 ( .A(sa22[7]), .B(sa22[6]), .Z(n5877) );
  HS65_LL_NOR2X6 U17794 ( .A(sa23[7]), .B(sa23[6]), .Z(n7460) );
  HS65_LL_NOR2X6 U17795 ( .A(sa00[7]), .B(sa00[6]), .Z(n5803) );
  HS65_LL_NOR2X6 U17796 ( .A(sa01[7]), .B(sa01[6]), .Z(n7395) );
  HS65_LL_NOR2X6 U17797 ( .A(sa20[1]), .B(sa20[0]), .Z(n9028) );
  HS65_LL_NOR2X6 U17798 ( .A(sa13[1]), .B(sa13[0]), .Z(n9086) );
  HS65_LL_NOR2X6 U17799 ( .A(sa11[5]), .B(sa11[4]), .Z(n5922) );
  HS65_LL_NOR2X6 U17800 ( .A(sa33[5]), .B(sa33[4]), .Z(n5740) );
  HS65_LL_NOR2X6 U17801 ( .A(sa12[5]), .B(sa12[4]), .Z(n7514) );
  HS65_LL_NOR2X6 U17802 ( .A(sa22[5]), .B(sa22[4]), .Z(n5863) );
  HS65_LL_NOR2X6 U17803 ( .A(sa23[5]), .B(sa23[4]), .Z(n7457) );
  HS65_LL_NOR2X6 U17804 ( .A(sa30[5]), .B(sa30[4]), .Z(n7332) );
  HS65_LL_NOR2X6 U17805 ( .A(sa00[5]), .B(sa00[4]), .Z(n5802) );
  HS65_LL_NOR2X6 U17806 ( .A(sa01[5]), .B(sa01[4]), .Z(n7394) );
  HS65_LL_NOR2X6 U17807 ( .A(w3[25]), .B(w3[24]), .Z(n2608) );
  HS65_LL_NOR2X6 U17808 ( .A(w3[17]), .B(w3[16]), .Z(n1480) );
  HS65_LL_NOR2X6 U17809 ( .A(w3[9]), .B(w3[8]), .Z(n1856) );
  HS65_LL_NOR2X6 U17810 ( .A(n899), .B(w3[27]), .Z(n2604) );
  HS65_LL_NOR2X6 U17811 ( .A(n858), .B(w3[19]), .Z(n1476) );
  HS65_LL_NOR2X6 U17812 ( .A(n776), .B(w3[3]), .Z(n2228) );
  HS65_LL_OAI22X6 U17813 ( .A(n2741), .B(n9136), .C(n9127), .D(n2742), .Z(N51)
         );
  HS65_LLS_XNOR2X6 U17814 ( .A(w3[9]), .B(text_in_r[9]), .Z(n2741) );
  HS65_LLS_XNOR3X2 U17815 ( .A(n2712), .B(n2743), .C(n2744), .Z(n2742) );
  HS65_LLS_XOR3X2 U17816 ( .A(n2663), .B(n816), .C(n183), .Z(n2743) );
  HS65_LL_NOR2X6 U17817 ( .A(w3[29]), .B(w3[28]), .Z(n2593) );
  HS65_LL_NOR2X6 U17818 ( .A(w3[13]), .B(w3[12]), .Z(n1841) );
  HS65_LL_NOR2X6 U17819 ( .A(w3[21]), .B(w3[20]), .Z(n1465) );
  HS65_LL_NOR2X6 U17820 ( .A(w3[5]), .B(w3[4]), .Z(n2217) );
  HS65_LL_OAI22X6 U17821 ( .A(n2667), .B(n9131), .C(n9128), .D(n2668), .Z(N83)
         );
  HS65_LLS_XNOR2X6 U17822 ( .A(w3[25]), .B(text_in_r[25]), .Z(n2667) );
  HS65_LLS_XNOR3X2 U17823 ( .A(n2669), .B(n2670), .C(n2671), .Z(n2668) );
  HS65_LLS_XOR3X2 U17824 ( .A(n2673), .B(w3[25]), .C(n2674), .Z(n2670) );
  HS65_LL_OAI22X6 U17825 ( .A(n5963), .B(n9130), .C(n9124), .D(n5964), .Z(N211) );
  HS65_LLS_XNOR2X6 U17826 ( .A(w1[25]), .B(text_in_r[89]), .Z(n5963) );
  HS65_LLS_XNOR3X2 U17827 ( .A(n5965), .B(n5966), .C(n5967), .Z(n5964) );
  HS65_LLS_XNOR2X6 U17828 ( .A(n3006), .B(n272), .Z(n5967) );
  HS65_LL_OAI22X6 U17829 ( .A(n4370), .B(n9135), .C(n9126), .D(n4371), .Z(N275) );
  HS65_LLS_XNOR2X6 U17830 ( .A(w0[25]), .B(text_in_r[121]), .Z(n4370) );
  HS65_LLS_XNOR3X2 U17831 ( .A(n4372), .B(n4373), .C(n4374), .Z(n4371) );
  HS65_LLS_XNOR2X6 U17832 ( .A(n3209), .B(n447), .Z(n4374) );
  HS65_LL_NOR2X6 U17833 ( .A(w3[15]), .B(w3[14]), .Z(n1834) );
  HS65_LL_NOR2X6 U17834 ( .A(n838), .B(w3[14]), .Z(n1840) );
  HS65_LL_NOR2X6 U17835 ( .A(w3[31]), .B(w3[30]), .Z(n2586) );
  HS65_LL_NOR2X6 U17836 ( .A(n920), .B(w3[30]), .Z(n2592) );
  HS65_LL_NOR2X6 U17837 ( .A(n817), .B(w3[11]), .Z(n1852) );
  HS65_LLS_XNOR2X6 U17838 ( .A(n2233), .B(w0[7]), .Z(n1001) );
  HS65_LL_NOR3X4 U17839 ( .A(n2234), .B(n2235), .C(n2236), .Z(n2233) );
  HS65_LL_NAND4ABX3 U17840 ( .A(n2247), .B(n2248), .C(n2249), .D(n2250), .Z(
        n2235) );
  HS65_LL_OAI212X5 U17841 ( .A(n2237), .B(n2238), .C(n2239), .D(n2240), .E(
        n2241), .Z(n2236) );
  HS65_LL_NOR2X6 U17842 ( .A(n271), .B(sa22[1]), .Z(n5872) );
  HS65_LL_NOR2X6 U17843 ( .A(n488), .B(sa11[1]), .Z(n5931) );
  HS65_LL_NOR2X6 U17844 ( .A(n49), .B(sa33[1]), .Z(n5746) );
  HS65_LL_NOR2X6 U17845 ( .A(n704), .B(sa00[1]), .Z(n5808) );
  HS65_LL_NOR2X6 U17846 ( .A(n313), .B(sa12[1]), .Z(n7523) );
  HS65_LL_NOR2X6 U17847 ( .A(n528), .B(sa01[1]), .Z(n7400) );
  HS65_LL_NOR2X6 U17848 ( .A(n571), .B(sa30[1]), .Z(n7338) );
  HS65_LL_NOR2X6 U17849 ( .A(n93), .B(sa23[1]), .Z(n7456) );
  HS65_LL_NOR2X6 U17850 ( .A(sa10[1]), .B(sa10[0]), .Z(n4284) );
  HS65_LL_NOR2X6 U17851 ( .A(n182), .B(sa03[0]), .Z(n4157) );
  HS65_LL_NOR2X6 U17852 ( .A(n619), .B(sa20[1]), .Z(n9041) );
  HS65_LL_NOR2X6 U17853 ( .A(n139), .B(sa13[1]), .Z(n9099) );
  HS65_LL_NOR2X6 U17854 ( .A(n27), .B(sa33[5]), .Z(n5738) );
  HS65_LL_NOR2X6 U17855 ( .A(n549), .B(sa30[5]), .Z(n7330) );
  HS65_LLS_XNOR2X6 U17856 ( .A(n1903), .B(w0[13]), .Z(n995) );
  HS65_LL_NOR3X4 U17857 ( .A(n1904), .B(n1905), .C(n1906), .Z(n1903) );
  HS65_LL_OAI212X5 U17858 ( .A(n1907), .B(n1908), .C(n1909), .D(n1862), .E(
        n1910), .Z(n1906) );
  HS65_LL_NAND4ABX3 U17859 ( .A(n1916), .B(n1917), .C(n1918), .D(n1919), .Z(
        n1905) );
  HS65_LLS_XNOR2X6 U17860 ( .A(n1945), .B(w0[12]), .Z(n996) );
  HS65_LL_NOR3X4 U17861 ( .A(n1946), .B(n1947), .C(n1948), .Z(n1945) );
  HS65_LL_OAI212X5 U17862 ( .A(n1949), .B(n1864), .C(n1950), .D(n1951), .E(
        n1952), .Z(n1948) );
  HS65_LL_NAND4ABX3 U17863 ( .A(n1953), .B(n1954), .C(n1955), .D(n1956), .Z(
        n1947) );
  HS65_LLS_XNOR2X6 U17864 ( .A(n1481), .B(w0[23]), .Z(n985) );
  HS65_LL_NOR3X4 U17865 ( .A(n1482), .B(n1483), .C(n1484), .Z(n1481) );
  HS65_LL_OAI212X5 U17866 ( .A(n1485), .B(n1486), .C(n1487), .D(n1488), .E(
        n1489), .Z(n1484) );
  HS65_LL_NAND4ABX3 U17867 ( .A(n1495), .B(n1496), .C(n1497), .D(n1498), .Z(
        n1483) );
  HS65_LLS_XNOR2X6 U17868 ( .A(n2502), .B(w0[2]), .Z(n1006) );
  HS65_LL_NOR4ABX2 U17869 ( .A(n2503), .B(n2504), .C(n2505), .D(n2506), .Z(
        n2502) );
  HS65_LL_CBI4I1X5 U17870 ( .A(n2291), .B(n2239), .C(n2273), .D(n2469), .Z(
        n2506) );
  HS65_LL_AOI212X4 U17871 ( .A(n893), .B(n912), .C(n901), .D(n2251), .E(n2521), 
        .Z(n2504) );
  HS65_LL_NOR2X6 U17872 ( .A(sa32[7]), .B(sa32[6]), .Z(n4217) );
  HS65_LL_NOR2X6 U17873 ( .A(n897), .B(w3[25]), .Z(n2603) );
  HS65_LL_NOR2X6 U17874 ( .A(sa20[3]), .B(sa20[2]), .Z(n9027) );
  HS65_LL_NOR2X6 U17875 ( .A(sa13[3]), .B(sa13[2]), .Z(n9085) );
  HS65_LL_NOR2X6 U17876 ( .A(sa03[5]), .B(sa03[4]), .Z(n4140) );
  HS65_LL_NOR2X6 U17877 ( .A(sa32[1]), .B(sa32[0]), .Z(n4209) );
  HS65_LL_NOR2X6 U17878 ( .A(sa21[1]), .B(sa21[0]), .Z(n4343) );
  HS65_LL_NOR2X6 U17879 ( .A(n159), .B(sa03[6]), .Z(n4151) );
  HS65_LL_NOR2X6 U17880 ( .A(n663), .B(sa10[3]), .Z(n4282) );
  HS65_LL_NOR2X6 U17881 ( .A(n138), .B(sa13[3]), .Z(n9098) );
  HS65_LL_NOR2X6 U17882 ( .A(n618), .B(sa20[3]), .Z(n9040) );
  HS65_LL_NOR2X6 U17883 ( .A(sa31[1]), .B(sa31[0]), .Z(n8971) );
  HS65_LL_NOR2X6 U17884 ( .A(n358), .B(sa02[0]), .Z(n8917) );
  HS65_LL_NOR2X6 U17885 ( .A(n270), .B(sa22[3]), .Z(n5851) );
  HS65_LL_NOR2X6 U17886 ( .A(n487), .B(sa11[3]), .Z(n5910) );
  HS65_LL_NOR2X6 U17887 ( .A(n92), .B(sa23[3]), .Z(n7443) );
  HS65_LL_NOR2X6 U17888 ( .A(n312), .B(sa12[3]), .Z(n7502) );
  HS65_LL_NOR2X6 U17889 ( .A(n703), .B(sa00[3]), .Z(n5804) );
  HS65_LL_NOR2X6 U17890 ( .A(n527), .B(sa01[3]), .Z(n7396) );
  HS65_LL_NOR2X6 U17891 ( .A(sa22[1]), .B(sa22[0]), .Z(n5870) );
  HS65_LL_NOR2X6 U17892 ( .A(sa11[1]), .B(sa11[0]), .Z(n5929) );
  HS65_LL_NOR2X6 U17893 ( .A(sa00[1]), .B(sa00[0]), .Z(n5805) );
  HS65_LL_NOR2X6 U17894 ( .A(sa23[1]), .B(sa23[0]), .Z(n7453) );
  HS65_LL_NOR2X6 U17895 ( .A(sa12[1]), .B(sa12[0]), .Z(n7521) );
  HS65_LL_NOR2X6 U17896 ( .A(sa01[1]), .B(sa01[0]), .Z(n7397) );
  HS65_LL_NOR2X6 U17897 ( .A(n338), .B(sa02[5]), .Z(n8908) );
  HS65_LL_NOR2X6 U17898 ( .A(sa33[7]), .B(sa33[6]), .Z(n5741) );
  HS65_LL_NOR2X6 U17899 ( .A(sa30[7]), .B(sa30[6]), .Z(n7333) );
  HS65_LL_NOR2X6 U17900 ( .A(n774), .B(w3[1]), .Z(n2227) );
  HS65_LL_NOR2X6 U17901 ( .A(n856), .B(w3[17]), .Z(n1475) );
  HS65_LLS_XNOR2X6 U17902 ( .A(w2[24]), .B(n1080), .Z(n1024) );
  HS65_LLS_XNOR2X6 U17903 ( .A(w2[5]), .B(n1099), .Z(n1062) );
  HS65_LLS_XNOR2X6 U17904 ( .A(w2[22]), .B(n1082), .Z(n1028) );
  HS65_LLS_XNOR2X6 U17905 ( .A(w2[10]), .B(n1094), .Z(n1052) );
  HS65_LLS_XNOR2X6 U17906 ( .A(w2[4]), .B(n1100), .Z(n1064) );
  HS65_LLS_XNOR2X6 U17907 ( .A(w2[12]), .B(n1092), .Z(n1048) );
  HS65_LLS_XNOR2X6 U17908 ( .A(w2[1]), .B(n1103), .Z(n1070) );
  HS65_LLS_XNOR2X6 U17909 ( .A(w2[15]), .B(n1089), .Z(n1042) );
  HS65_LLS_XNOR2X6 U17910 ( .A(w0[0]), .B(n2549), .Z(n1008) );
  HS65_LL_NAND4ABX3 U17911 ( .A(n2550), .B(n2551), .C(n2552), .D(n2553), .Z(
        n2549) );
  HS65_LL_MX41X7 U17912 ( .D0(n893), .S0(n910), .D1(n894), .S1(n902), .D2(n913), .S2(n886), .D3(n914), .S3(n2313), .Z(n2551) );
  HS65_LL_NOR4ABX2 U17913 ( .A(n2311), .B(n2446), .C(n2554), .D(n2460), .Z(
        n2553) );
  HS65_LLS_XNOR2X6 U17914 ( .A(w0[8]), .B(n2173), .Z(n1000) );
  HS65_LL_NAND4ABX3 U17915 ( .A(n2174), .B(n2175), .C(n2176), .D(n2177), .Z(
        n2173) );
  HS65_LL_MX41X7 U17916 ( .D0(n770), .S0(n787), .D1(n771), .S1(n779), .D2(n790), .S2(n763), .D3(n791), .S3(n1937), .Z(n2175) );
  HS65_LL_NOR4ABX2 U17917 ( .A(n1935), .B(n2070), .C(n2178), .D(n2084), .Z(
        n2177) );
  HS65_LLS_XNOR2X6 U17918 ( .A(w2[8]), .B(n1096), .Z(n1056) );
  HS65_LL_NOR2X6 U17919 ( .A(n815), .B(w3[9]), .Z(n1851) );
  HS65_LL_IVX9 U17920 ( .A(w3[14]), .Z(n837) );
  HS65_LL_IVX9 U17921 ( .A(w3[30]), .Z(n919) );
  HS65_LL_IVX9 U17922 ( .A(w3[10]), .Z(n817) );
  HS65_LL_IVX9 U17923 ( .A(w3[29]), .Z(n918) );
  HS65_LL_IVX9 U17924 ( .A(w3[13]), .Z(n836) );
  HS65_LLS_XNOR2X6 U17925 ( .A(w0[9]), .B(n2148), .Z(n999) );
  HS65_LL_NAND4ABX3 U17926 ( .A(n2149), .B(n2150), .C(n2151), .D(n2152), .Z(
        n2148) );
  HS65_LL_CB4I6X9 U17927 ( .A(n762), .B(n767), .C(n789), .D(n2086), .Z(n2149)
         );
  HS65_LL_AOI222X2 U17928 ( .A(n781), .B(n759), .C(n778), .D(n2171), .E(n790), 
        .F(n758), .Z(n2151) );
  HS65_LLS_XNOR2X6 U17929 ( .A(w2[31]), .B(n1073), .Z(n1010) );
  HS65_LLS_XNOR2X6 U17930 ( .A(w2[13]), .B(n1091), .Z(n1046) );
  HS65_LLS_XNOR2X6 U17931 ( .A(w2[29]), .B(n1075), .Z(n1014) );
  HS65_LLS_XNOR2X6 U17932 ( .A(w2[14]), .B(n1090), .Z(n1044) );
  HS65_LLS_XNOR2X6 U17933 ( .A(w2[3]), .B(n1101), .Z(n1066) );
  HS65_LL_IVX9 U17934 ( .A(w3[11]), .Z(n818) );
  HS65_LL_IVX9 U17935 ( .A(w3[9]), .Z(n816) );
  HS65_LLS_XNOR2X6 U17936 ( .A(w0[11]), .B(n2007), .Z(n997) );
  HS65_LL_NAND4ABX3 U17937 ( .A(n2008), .B(n2009), .C(n2010), .D(n2011), .Z(
        n2007) );
  HS65_LL_AOI212X4 U17938 ( .A(n773), .B(n2012), .C(n789), .D(n1989), .E(n2013), .Z(n2011) );
  HS65_LL_MX41X7 U17939 ( .D0(n760), .S0(n784), .D1(n788), .S1(n772), .D2(n758), .S2(n779), .D3(n790), .S3(n1937), .Z(n2009) );
  HS65_LLS_XNOR2X6 U17940 ( .A(w2[25]), .B(n1079), .Z(n1022) );
  HS65_LLS_XNOR2X6 U17941 ( .A(w2[9]), .B(n1095), .Z(n1054) );
  HS65_LLS_XNOR2X6 U17942 ( .A(w2[11]), .B(n1093), .Z(n1050) );
  HS65_LLS_XNOR2X6 U17943 ( .A(w0[22]), .B(n1508), .Z(n986) );
  HS65_LL_NAND4ABX3 U17944 ( .A(n1509), .B(n1510), .C(n1511), .D(n1512), .Z(
        n1508) );
  HS65_LL_AOI212X4 U17945 ( .A(n832), .B(n798), .C(n829), .D(n810), .E(n1518), 
        .Z(n1511) );
  HS65_LL_CBI4I1X5 U17946 ( .A(n1524), .B(n1486), .C(n1525), .D(n1526), .Z(
        n1509) );
  HS65_LLS_XNOR2X6 U17947 ( .A(w2[0]), .B(n1104), .Z(n1072) );
  HS65_LLS_XNOR2X6 U17948 ( .A(w2[23]), .B(n1081), .Z(n1026) );
  HS65_LLS_XNOR2X6 U17949 ( .A(w2[2]), .B(n1102), .Z(n1068) );
  HS65_LLS_XNOR2X6 U17950 ( .A(w2[6]), .B(n1098), .Z(n1060) );
  HS65_LLS_XNOR2X6 U17951 ( .A(w2[27]), .B(n1077), .Z(n1018) );
  HS65_LLS_XNOR2X6 U17952 ( .A(w2[17]), .B(n1087), .Z(n1038) );
  HS65_LLS_XNOR2X6 U17953 ( .A(w2[19]), .B(n1085), .Z(n1034) );
  HS65_LLS_XNOR2X6 U17954 ( .A(w2[20]), .B(n1084), .Z(n1032) );
  HS65_LLS_XNOR2X6 U17955 ( .A(w2[16]), .B(n1088), .Z(n1040) );
  HS65_LLS_XNOR2X6 U17956 ( .A(w2[7]), .B(n1097), .Z(n1058) );
  HS65_LLS_XNOR2X6 U17957 ( .A(w2[18]), .B(n1086), .Z(n1036) );
  HS65_LLS_XNOR2X6 U17958 ( .A(w2[21]), .B(n1083), .Z(n1030) );
  HS65_LL_NOR2X6 U17959 ( .A(n70), .B(sa23[7]), .Z(n7468) );
  HS65_LL_NOR2X6 U17960 ( .A(n248), .B(sa22[7]), .Z(n5875) );
  HS65_LL_NOR2X6 U17961 ( .A(n465), .B(sa11[7]), .Z(n5934) );
  HS65_LL_NOR2X6 U17962 ( .A(n290), .B(sa12[7]), .Z(n7526) );
  HS65_LL_NOR2X6 U17963 ( .A(n505), .B(sa01[7]), .Z(n7399) );
  HS65_LL_NOR2X6 U17964 ( .A(n681), .B(sa00[7]), .Z(n5807) );
  HS65_LL_IVX9 U17965 ( .A(w3[26]), .Z(n899) );
  HS65_LL_IVX9 U17966 ( .A(w3[31]), .Z(n920) );
  HS65_LL_IVX9 U17967 ( .A(w3[28]), .Z(n917) );
  HS65_LL_IVX9 U17968 ( .A(w3[12]), .Z(n835) );
  HS65_LL_IVX9 U17969 ( .A(w3[16]), .Z(n856) );
  HS65_LL_IVX9 U17970 ( .A(w3[24]), .Z(n897) );
  HS65_LL_IVX9 U17971 ( .A(w3[8]), .Z(n815) );
  HS65_LL_IVX9 U17972 ( .A(w3[20]), .Z(n876) );
  HS65_LL_IVX9 U17973 ( .A(w3[4]), .Z(n794) );
  HS65_LL_IVX9 U17974 ( .A(w3[27]), .Z(n900) );
  HS65_LL_IVX9 U17975 ( .A(w3[1]), .Z(n775) );
  HS65_LLS_XNOR2X6 U17976 ( .A(w1[3]), .B(n1005), .Z(n1101) );
  HS65_LLS_XNOR2X6 U17977 ( .A(w1[27]), .B(n981), .Z(n1077) );
  HS65_LL_IVX9 U17978 ( .A(w3[19]), .Z(n859) );
  HS65_LL_IVX9 U17979 ( .A(w3[3]), .Z(n777) );
  HS65_LL_IVX9 U17980 ( .A(w3[17]), .Z(n857) );
  HS65_LL_IVX9 U17981 ( .A(w3[7]), .Z(n797) );
  HS65_LL_IVX9 U17982 ( .A(w3[23]), .Z(n879) );
  HS65_LLS_XNOR2X6 U17983 ( .A(w1[17]), .B(n991), .Z(n1087) );
  HS65_LLS_XNOR2X6 U17984 ( .A(w1[19]), .B(n989), .Z(n1085) );
  HS65_LLS_XNOR2X6 U17985 ( .A(w1[16]), .B(n992), .Z(n1088) );
  HS65_LLS_XNOR2X6 U17986 ( .A(w1[24]), .B(n984), .Z(n1080) );
  HS65_LLS_XOR2X6 U17987 ( .A(n995), .B(w1[13]), .Z(n1091) );
  HS65_LLS_XOR2X6 U17988 ( .A(n979), .B(w1[29]), .Z(n1075) );
  HS65_LLS_XOR2X6 U17989 ( .A(n1001), .B(w1[7]), .Z(n1097) );
  HS65_LLS_XNOR2X6 U17990 ( .A(w2[26]), .B(n1078), .Z(n1020) );
  HS65_LLS_XNOR2X6 U17991 ( .A(w2[30]), .B(n1074), .Z(n1012) );
  HS65_LLS_XNOR2X6 U17992 ( .A(w2[28]), .B(n1076), .Z(n1016) );
  HS65_LL_NOR2X6 U17993 ( .A(n48), .B(sa33[3]), .Z(n5742) );
  HS65_LL_NOR2X6 U17994 ( .A(n570), .B(sa30[3]), .Z(n7334) );
  HS65_LL_IVX9 U17995 ( .A(w3[0]), .Z(n774) );
  HS65_LL_IVX9 U17996 ( .A(w3[22]), .Z(n878) );
  HS65_LL_IVX9 U17997 ( .A(w3[6]), .Z(n796) );
  HS65_LL_IVX9 U17998 ( .A(w3[2]), .Z(n776) );
  HS65_LL_IVX9 U17999 ( .A(w3[18]), .Z(n858) );
  HS65_LL_IVX9 U18000 ( .A(w3[15]), .Z(n838) );
  HS65_LL_IVX9 U18001 ( .A(w3[25]), .Z(n898) );
  HS65_LLS_XNOR2X6 U18002 ( .A(w1[9]), .B(n999), .Z(n1095) );
  HS65_LLS_XNOR2X6 U18003 ( .A(w1[14]), .B(n994), .Z(n1090) );
  HS65_LLS_XNOR2X6 U18004 ( .A(w1[1]), .B(n1007), .Z(n1103) );
  HS65_LL_IVX9 U18005 ( .A(w3[21]), .Z(n877) );
  HS65_LL_IVX9 U18006 ( .A(w3[5]), .Z(n795) );
  HS65_LLS_XNOR2X6 U18007 ( .A(w1[11]), .B(n997), .Z(n1093) );
  HS65_LLS_XNOR2X6 U18008 ( .A(w1[0]), .B(n1008), .Z(n1104) );
  HS65_LLS_XNOR2X6 U18009 ( .A(w1[8]), .B(n1000), .Z(n1096) );
  HS65_LLS_XNOR2X6 U18010 ( .A(w1[6]), .B(n1002), .Z(n1098) );
  HS65_LLS_XNOR2X6 U18011 ( .A(w1[22]), .B(n986), .Z(n1082) );
  HS65_LL_NOR2X6 U18012 ( .A(n446), .B(sa21[1]), .Z(n4338) );
  HS65_LL_NOR2X6 U18013 ( .A(n228), .B(sa32[1]), .Z(n4214) );
  HS65_LLS_XOR2X6 U18014 ( .A(n1004), .B(w1[4]), .Z(n1100) );
  HS65_LLS_XOR2X6 U18015 ( .A(n996), .B(w1[12]), .Z(n1092) );
  HS65_LLS_XOR2X6 U18016 ( .A(n985), .B(w1[23]), .Z(n1081) );
  HS65_LLS_XOR2X6 U18017 ( .A(n1006), .B(w1[2]), .Z(n1102) );
  HS65_LLS_XOR2X6 U18018 ( .A(n980), .B(w1[28]), .Z(n1076) );
  HS65_LLS_XOR2X6 U18019 ( .A(n988), .B(w1[20]), .Z(n1084) );
  HS65_LLS_XOR2X6 U18020 ( .A(n990), .B(w1[18]), .Z(n1086) );
  HS65_LLS_XOR2X6 U18021 ( .A(n987), .B(w1[21]), .Z(n1083) );
  HS65_LLS_XOR2X6 U18022 ( .A(n1003), .B(w1[5]), .Z(n1099) );
  HS65_LL_AO22X9 U18023 ( .A(key[28]), .B(n9140), .C(n1015), .D(n9118), .Z(
        \u0/N268 ) );
  HS65_LLS_XNOR2X6 U18024 ( .A(w3[28]), .B(n1016), .Z(n1015) );
  HS65_LL_AO22X9 U18025 ( .A(key[4]), .B(n9137), .C(n1063), .D(n9146), .Z(
        \u0/N244 ) );
  HS65_LLS_XNOR2X6 U18026 ( .A(w3[4]), .B(n1064), .Z(n1063) );
  HS65_LL_AO22X9 U18027 ( .A(key[26]), .B(n9140), .C(n1019), .D(n9144), .Z(
        \u0/N266 ) );
  HS65_LLS_XNOR2X6 U18028 ( .A(w3[26]), .B(n1020), .Z(n1019) );
  HS65_LL_AO22X9 U18029 ( .A(key[27]), .B(n9140), .C(n1017), .D(n9148), .Z(
        \u0/N267 ) );
  HS65_LLS_XNOR2X6 U18030 ( .A(w3[27]), .B(n1018), .Z(n1017) );
  HS65_LLS_XOR2X6 U18031 ( .A(n977), .B(w1[31]), .Z(n1073) );
  HS65_LLS_XOR2X6 U18032 ( .A(n998), .B(w1[10]), .Z(n1094) );
  HS65_LLS_XOR2X6 U18033 ( .A(n993), .B(w1[15]), .Z(n1089) );
  HS65_LLS_XOR2X6 U18034 ( .A(n982), .B(w1[26]), .Z(n1078) );
  HS65_LL_AND2X4 U18035 ( .A(sa22[7]), .B(sa22[6]), .Z(n5855) );
  HS65_LL_AND2X4 U18036 ( .A(sa11[7]), .B(sa11[6]), .Z(n5914) );
  HS65_LL_AND2X4 U18037 ( .A(sa33[7]), .B(sa33[6]), .Z(n5739) );
  HS65_LL_AND2X4 U18038 ( .A(sa12[7]), .B(sa12[6]), .Z(n7506) );
  HS65_LL_AND2X4 U18039 ( .A(sa30[7]), .B(sa30[6]), .Z(n7331) );
  HS65_LL_AND2X4 U18040 ( .A(sa01[7]), .B(sa01[6]), .Z(n7393) );
  HS65_LL_AND2X4 U18041 ( .A(sa23[7]), .B(sa23[6]), .Z(n7447) );
  HS65_LL_AO22X9 U18042 ( .A(key[29]), .B(n9140), .C(n1013), .D(n9146), .Z(
        \u0/N269 ) );
  HS65_LLS_XNOR2X6 U18043 ( .A(w3[29]), .B(n1014), .Z(n1013) );
  HS65_LL_AO22X9 U18044 ( .A(key[11]), .B(n9137), .C(n1049), .D(n9146), .Z(
        \u0/N251 ) );
  HS65_LLS_XNOR2X6 U18045 ( .A(w3[11]), .B(n1050), .Z(n1049) );
  HS65_LL_AO22X9 U18046 ( .A(key[9]), .B(n9137), .C(n1053), .D(n9146), .Z(
        \u0/N249 ) );
  HS65_LLS_XNOR2X6 U18047 ( .A(w3[9]), .B(n1054), .Z(n1053) );
  HS65_LL_AND2X4 U18048 ( .A(sa33[5]), .B(sa33[4]), .Z(n5744) );
  HS65_LL_AND2X4 U18049 ( .A(sa30[5]), .B(sa30[4]), .Z(n7336) );
  HS65_LL_AND2X4 U18050 ( .A(sa33[5]), .B(n27), .Z(n5752) );
  HS65_LL_AND2X4 U18051 ( .A(sa30[5]), .B(n549), .Z(n7344) );
  HS65_LL_AND2X4 U18052 ( .A(sa11[5]), .B(sa11[4]), .Z(n5924) );
  HS65_LL_AND2X4 U18053 ( .A(sa22[5]), .B(sa22[4]), .Z(n5865) );
  HS65_LL_AND2X4 U18054 ( .A(sa12[5]), .B(sa12[4]), .Z(n7516) );
  HS65_LL_AND2X4 U18055 ( .A(sa23[5]), .B(sa23[4]), .Z(n7459) );
  HS65_LL_AND2X4 U18056 ( .A(sa01[5]), .B(sa01[4]), .Z(n7398) );
  HS65_LL_AND2X4 U18057 ( .A(sa00[5]), .B(sa00[4]), .Z(n5806) );
  HS65_LL_AND2X4 U18058 ( .A(sa22[1]), .B(sa22[0]), .Z(n5852) );
  HS65_LL_AND2X4 U18059 ( .A(sa11[1]), .B(sa11[0]), .Z(n5911) );
  HS65_LL_AND2X4 U18060 ( .A(sa23[1]), .B(sa23[0]), .Z(n7444) );
  HS65_LL_AND2X4 U18061 ( .A(sa12[1]), .B(sa12[0]), .Z(n7503) );
  HS65_LL_AND2X4 U18062 ( .A(sa01[1]), .B(sa01[0]), .Z(n7382) );
  HS65_LL_AND2X4 U18063 ( .A(sa00[1]), .B(sa00[0]), .Z(n5790) );
  HS65_LL_AND2X4 U18064 ( .A(sa10[0]), .B(sa10[1]), .Z(n4272) );
  HS65_LL_OAI22X6 U18065 ( .A(n2899), .B(n9136), .C(n9127), .D(n2900), .Z(N40)
         );
  HS65_LLS_XNOR2X6 U18066 ( .A(w3[6]), .B(text_in_r[6]), .Z(n2899) );
  HS65_LLS_XOR3X2 U18067 ( .A(n2636), .B(n2690), .C(n2901), .Z(n2900) );
  HS65_LLS_XNOR2X6 U18068 ( .A(w3[6]), .B(n2631), .Z(n2901) );
  HS65_LL_OAI22X6 U18069 ( .A(n2683), .B(n9131), .C(n9128), .D(n2684), .Z(N72)
         );
  HS65_LLS_XNOR2X6 U18070 ( .A(w3[22]), .B(text_in_r[22]), .Z(n2683) );
  HS65_LLS_XOR3X2 U18071 ( .A(n2643), .B(n2685), .C(n2686), .Z(n2684) );
  HS65_LLS_XNOR2X6 U18072 ( .A(w3[22]), .B(n2687), .Z(n2686) );
  HS65_LL_OAI22X6 U18073 ( .A(n2704), .B(n9131), .C(n9128), .D(n2705), .Z(N68)
         );
  HS65_LLS_XNOR2X6 U18074 ( .A(w3[18]), .B(text_in_r[18]), .Z(n2704) );
  HS65_LLS_XOR3X2 U18075 ( .A(n2669), .B(n2706), .C(n2707), .Z(n2705) );
  HS65_LLS_XNOR2X6 U18076 ( .A(w3[18]), .B(n2708), .Z(n2707) );
  HS65_LL_OAI22X6 U18077 ( .A(n3899), .B(n9136), .C(n9127), .D(n3900), .Z(N36)
         );
  HS65_LLS_XNOR2X6 U18078 ( .A(w3[2]), .B(text_in_r[2]), .Z(n3899) );
  HS65_LLS_XOR3X2 U18079 ( .A(n2665), .B(n2712), .C(n3901), .Z(n3900) );
  HS65_LLS_XNOR2X6 U18080 ( .A(w3[2]), .B(n141), .Z(n3901) );
  HS65_LL_IVX9 U18081 ( .A(sa10[6]), .Z(n641) );
  HS65_LL_IVX9 U18082 ( .A(sa02[6]), .Z(n336) );
  HS65_LL_IVX9 U18083 ( .A(sa32[6]), .Z(n205) );
  HS65_LL_IVX9 U18084 ( .A(sa03[6]), .Z(n160) );
  HS65_LL_IVX9 U18085 ( .A(sa20[4]), .Z(n597) );
  HS65_LL_IVX9 U18086 ( .A(sa31[6]), .Z(n380) );
  HS65_LL_IVX9 U18087 ( .A(sa13[4]), .Z(n117) );
  HS65_LL_IVX9 U18088 ( .A(sa02[0]), .Z(n359) );
  HS65_LL_IVX9 U18089 ( .A(sa13[2]), .Z(n138) );
  HS65_LL_IVX9 U18090 ( .A(sa20[2]), .Z(n618) );
  HS65_LL_IVX9 U18091 ( .A(sa22[2]), .Z(n270) );
  HS65_LL_IVX9 U18092 ( .A(sa11[2]), .Z(n487) );
  HS65_LL_IVX9 U18093 ( .A(sa33[2]), .Z(n48) );
  HS65_LL_IVX9 U18094 ( .A(sa00[2]), .Z(n703) );
  HS65_LL_IVX9 U18095 ( .A(sa21[0]), .Z(n446) );
  HS65_LL_IVX9 U18096 ( .A(sa10[2]), .Z(n663) );
  HS65_LL_IVX9 U18097 ( .A(sa32[0]), .Z(n228) );
  HS65_LL_IVX9 U18098 ( .A(sa03[4]), .Z(n162) );
  HS65_LL_IVX9 U18099 ( .A(sa02[4]), .Z(n338) );
  HS65_LL_IVX9 U18100 ( .A(sa31[4]), .Z(n382) );
  HS65_LL_IVX9 U18101 ( .A(sa12[2]), .Z(n312) );
  HS65_LL_IVX9 U18102 ( .A(sa01[2]), .Z(n527) );
  HS65_LL_IVX9 U18103 ( .A(sa30[2]), .Z(n570) );
  HS65_LL_IVX9 U18104 ( .A(sa23[2]), .Z(n92) );
  HS65_LL_IVX9 U18105 ( .A(sa31[0]), .Z(n403) );
  HS65_LL_IVX9 U18106 ( .A(sa21[6]), .Z(n423) );
  HS65_LL_IVX9 U18107 ( .A(sa32[5]), .Z(n206) );
  HS65_LL_IVX9 U18108 ( .A(sa21[5]), .Z(n424) );
  HS65_LL_IVX9 U18109 ( .A(sa10[5]), .Z(n642) );
  HS65_LL_IVX9 U18110 ( .A(sa03[3]), .Z(n176) );
  HS65_LL_IVX9 U18111 ( .A(sa13[7]), .Z(n114) );
  HS65_LL_IVX9 U18112 ( .A(sa20[7]), .Z(n594) );
  HS65_LL_OAI22X6 U18113 ( .A(n2729), .B(n9131), .C(n9127), .D(n2730), .Z(N54)
         );
  HS65_LLS_XNOR2X6 U18114 ( .A(w3[12]), .B(text_in_r[12]), .Z(n2729) );
  HS65_LLS_XOR3X2 U18115 ( .A(n2731), .B(n2697), .C(n2732), .Z(n2730) );
  HS65_LLS_XOR3X2 U18116 ( .A(w3[12]), .B(n2641), .C(n184), .Z(n2732) );
  HS65_LL_OAI22X6 U18117 ( .A(n2646), .B(n9131), .C(n9127), .D(n2647), .Z(N86)
         );
  HS65_LLS_XNOR2X6 U18118 ( .A(w3[28]), .B(text_in_r[28]), .Z(n2646) );
  HS65_LLS_XOR3X2 U18119 ( .A(n2648), .B(n2649), .C(n2650), .Z(n2647) );
  HS65_LLS_XOR3X2 U18120 ( .A(w3[28]), .B(n2651), .C(n2652), .Z(n2650) );
  HS65_LL_OAI22X6 U18121 ( .A(n2714), .B(n9131), .C(n9128), .D(n2715), .Z(N66)
         );
  HS65_LLS_XNOR2X6 U18122 ( .A(w3[16]), .B(text_in_r[16]), .Z(n2714) );
  HS65_LLS_XOR3X2 U18123 ( .A(n2695), .B(n2716), .C(n2717), .Z(n2715) );
  HS65_LLS_XNOR2X6 U18124 ( .A(w3[16]), .B(n2718), .Z(n2717) );
  HS65_LL_OAI22X6 U18125 ( .A(n2661), .B(n9131), .C(n9128), .D(n2662), .Z(N84)
         );
  HS65_LLS_XNOR2X6 U18126 ( .A(w3[26]), .B(text_in_r[26]), .Z(n2661) );
  HS65_LLS_XOR3X2 U18127 ( .A(n2663), .B(n2664), .C(n2665), .Z(n2662) );
  HS65_LLS_XOR3X2 U18128 ( .A(n2666), .B(n899), .C(n140), .Z(n2664) );
  HS65_LL_OAI22X6 U18129 ( .A(n2655), .B(n9131), .C(n9127), .D(n2656), .Z(N85)
         );
  HS65_LLS_XNOR2X6 U18130 ( .A(w3[27]), .B(text_in_r[27]), .Z(n2655) );
  HS65_LLS_XOR2X6 U18131 ( .A(n2657), .B(n2658), .Z(n2656) );
  HS65_LLS_XOR3X2 U18132 ( .A(w3[27]), .B(n141), .C(n184), .Z(n2657) );
  HS65_LL_AND2X4 U18133 ( .A(sa11[7]), .B(n465), .Z(n5923) );
  HS65_LL_AND2X4 U18134 ( .A(sa00[7]), .B(n681), .Z(n5810) );
  HS65_LL_AND2X4 U18135 ( .A(sa33[7]), .B(n26), .Z(n5748) );
  HS65_LL_AND2X4 U18136 ( .A(sa22[7]), .B(n248), .Z(n5864) );
  HS65_LL_AND2X4 U18137 ( .A(sa12[7]), .B(n290), .Z(n7515) );
  HS65_LL_AND2X4 U18138 ( .A(sa23[7]), .B(n70), .Z(n7458) );
  HS65_LL_AND2X4 U18139 ( .A(sa01[7]), .B(n505), .Z(n7402) );
  HS65_LL_AND2X4 U18140 ( .A(sa30[7]), .B(n548), .Z(n7340) );
  HS65_LL_IVX9 U18141 ( .A(sa21[4]), .Z(n425) );
  HS65_LL_IVX9 U18142 ( .A(sa13[6]), .Z(n115) );
  HS65_LL_IVX9 U18143 ( .A(sa20[6]), .Z(n595) );
  HS65_LL_IVX9 U18144 ( .A(sa32[4]), .Z(n207) );
  HS65_LL_IVX9 U18145 ( .A(sa10[4]), .Z(n643) );
  HS65_LL_IVX9 U18146 ( .A(sa03[2]), .Z(n181) );
  HS65_LL_AND2X4 U18147 ( .A(sa22[5]), .B(n249), .Z(n5876) );
  HS65_LL_AND2X4 U18148 ( .A(sa11[5]), .B(n466), .Z(n5935) );
  HS65_LL_AND2X4 U18149 ( .A(sa00[5]), .B(n682), .Z(n5814) );
  HS65_LL_AND2X4 U18150 ( .A(sa12[5]), .B(n291), .Z(n7527) );
  HS65_LL_AND2X4 U18151 ( .A(sa01[5]), .B(n506), .Z(n7406) );
  HS65_LL_AND2X4 U18152 ( .A(sa23[5]), .B(n71), .Z(n7469) );
  HS65_LL_IVX9 U18153 ( .A(sa10[3]), .Z(n662) );
  HS65_LL_IVX9 U18154 ( .A(sa10[7]), .Z(n632) );
  HS65_LL_IVX9 U18155 ( .A(sa13[5]), .Z(n116) );
  HS65_LL_IVX9 U18156 ( .A(sa20[5]), .Z(n596) );
  HS65_LL_IVX9 U18157 ( .A(sa02[5]), .Z(n337) );
  HS65_LL_IVX9 U18158 ( .A(sa31[7]), .Z(n379) );
  HS65_LL_IVX9 U18159 ( .A(sa31[5]), .Z(n381) );
  HS65_LL_IVX9 U18160 ( .A(sa02[1]), .Z(n358) );
  HS65_LL_IVX9 U18161 ( .A(sa13[3]), .Z(n133) );
  HS65_LL_IVX9 U18162 ( .A(sa22[3]), .Z(n269) );
  HS65_LL_IVX9 U18163 ( .A(sa11[3]), .Z(n486) );
  HS65_LL_IVX9 U18164 ( .A(sa33[3]), .Z(n43) );
  HS65_LL_IVX9 U18165 ( .A(sa00[3]), .Z(n698) );
  HS65_LL_IVX9 U18166 ( .A(sa21[7]), .Z(n414) );
  HS65_LL_IVX9 U18167 ( .A(sa21[1]), .Z(n445) );
  HS65_LL_IVX9 U18168 ( .A(sa32[7]), .Z(n204) );
  HS65_LL_IVX9 U18169 ( .A(sa03[5]), .Z(n161) );
  HS65_LL_IVX9 U18170 ( .A(sa03[7]), .Z(n159) );
  HS65_LL_IVX9 U18171 ( .A(sa20[3]), .Z(n613) );
  HS65_LL_IVX9 U18172 ( .A(sa02[7]), .Z(n331) );
  HS65_LL_IVX9 U18173 ( .A(sa12[3]), .Z(n311) );
  HS65_LL_IVX9 U18174 ( .A(sa01[3]), .Z(n522) );
  HS65_LL_IVX9 U18175 ( .A(sa30[3]), .Z(n565) );
  HS65_LL_IVX9 U18176 ( .A(sa23[3]), .Z(n87) );
  HS65_LL_IVX9 U18177 ( .A(sa31[1]), .Z(n402) );
  HS65_LL_IVX9 U18178 ( .A(sa32[1]), .Z(n227) );
  HS65_LL_OAI22X6 U18179 ( .A(n2738), .B(n9136), .C(n9127), .D(n2739), .Z(N52)
         );
  HS65_LLS_XNOR2X6 U18180 ( .A(w3[10]), .B(text_in_r[10]), .Z(n2738) );
  HS65_LLS_XNOR3X2 U18181 ( .A(n2713), .B(n2740), .C(n2706), .Z(n2739) );
  HS65_LLS_XOR3X2 U18182 ( .A(n2659), .B(n817), .C(n2673), .Z(n2740) );
  HS65_LL_OAI22X6 U18183 ( .A(n2734), .B(n9131), .C(n9127), .D(n2735), .Z(N53)
         );
  HS65_LLS_XNOR2X6 U18184 ( .A(w3[11]), .B(text_in_r[11]), .Z(n2734) );
  HS65_LLS_XOR2X6 U18185 ( .A(n2736), .B(n2737), .Z(n2735) );
  HS65_LLS_XOR3X2 U18186 ( .A(n2653), .B(n818), .C(n2708), .Z(n2736) );
  HS65_LL_OAI22X6 U18187 ( .A(n7566), .B(n9132), .C(n9126), .D(n7567), .Z(N136) );
  HS65_LLS_XNOR2X6 U18188 ( .A(w2[22]), .B(text_in_r[54]), .Z(n7566) );
  HS65_LLS_XOR3X2 U18189 ( .A(n7540), .B(n7568), .C(n7569), .Z(n7567) );
  HS65_LLS_XOR2X6 U18190 ( .A(w2[22]), .B(n2780), .Z(n7569) );
  HS65_LL_OAI22X6 U18191 ( .A(n7560), .B(n9132), .C(n9125), .D(n7561), .Z(N146) );
  HS65_LLS_XNOR2X6 U18192 ( .A(w2[24]), .B(text_in_r[56]), .Z(n7560) );
  HS65_LLS_XOR3X2 U18193 ( .A(n2623), .B(n7546), .C(n7562), .Z(n7561) );
  HS65_LLS_XOR2X6 U18194 ( .A(w2[24]), .B(n2750), .Z(n7562) );
  HS65_LL_OAI22X6 U18195 ( .A(n5954), .B(n9130), .C(n9124), .D(n5955), .Z(N213) );
  HS65_LLS_XNOR2X6 U18196 ( .A(w1[27]), .B(text_in_r[91]), .Z(n5954) );
  HS65_LLS_XOR3X2 U18197 ( .A(n5956), .B(n5957), .C(n5958), .Z(n5955) );
  HS65_LLS_XNOR3X2 U18198 ( .A(w1[27]), .B(n2761), .C(n2808), .Z(n5958) );
  HS65_LL_OAI22X6 U18199 ( .A(n8188), .B(n9132), .C(n9127), .D(n8189), .Z(N102) );
  HS65_LLS_XNOR2X6 U18200 ( .A(w2[4]), .B(text_in_r[36]), .Z(n8188) );
  HS65_LLS_XOR3X2 U18201 ( .A(n7544), .B(n8190), .C(n7582), .Z(n8189) );
  HS65_LLS_XNOR3X2 U18202 ( .A(w2[4]), .B(n2616), .C(n3002), .Z(n8190) );
  HS65_LL_OAI22X6 U18203 ( .A(n6707), .B(n9129), .C(n9122), .D(n6708), .Z(N165) );
  HS65_LLS_XNOR2X6 U18204 ( .A(w1[3]), .B(text_in_r[67]), .Z(n6707) );
  HS65_LLS_XOR3X2 U18205 ( .A(n5995), .B(n6709), .C(n6396), .Z(n6708) );
  HS65_LLS_XNOR3X2 U18206 ( .A(w1[3]), .B(n5957), .C(n3009), .Z(n6709) );
  HS65_LL_OAI22X6 U18207 ( .A(n6393), .B(n9129), .C(n9122), .D(n6394), .Z(N166) );
  HS65_LLS_XNOR2X6 U18208 ( .A(w1[4]), .B(text_in_r[68]), .Z(n6393) );
  HS65_LLS_XOR3X2 U18209 ( .A(n5992), .B(n6395), .C(n6396), .Z(n6394) );
  HS65_LLS_XNOR3X2 U18210 ( .A(w1[4]), .B(n5952), .C(n3205), .Z(n6395) );
  HS65_LL_OAI22X6 U18211 ( .A(n6014), .B(n9129), .C(n9123), .D(n6015), .Z(N182) );
  HS65_LLS_XNOR2X6 U18212 ( .A(w1[12]), .B(text_in_r[76]), .Z(n6014) );
  HS65_LLS_XOR3X2 U18213 ( .A(n6016), .B(n5988), .C(n6017), .Z(n6015) );
  HS65_LLS_XOR3X2 U18214 ( .A(w1[12]), .B(n2761), .C(n2785), .Z(n6017) );
  HS65_LL_OAI22X6 U18215 ( .A(n7594), .B(n9132), .C(n9126), .D(n7595), .Z(N121) );
  HS65_LLS_XNOR2X6 U18216 ( .A(w2[15]), .B(text_in_r[47]), .Z(n7594) );
  HS65_LLS_XOR3X2 U18217 ( .A(n2780), .B(n7596), .C(n7546), .Z(n7595) );
  HS65_LLS_XNOR3X2 U18218 ( .A(n2757), .B(w2[15]), .C(n2756), .Z(n7596) );
  HS65_LL_OAI22X6 U18219 ( .A(n4436), .B(n9135), .C(n9125), .D(n4437), .Z(N242) );
  HS65_LLS_XNOR2X6 U18220 ( .A(w0[8]), .B(text_in_r[104]), .Z(n4436) );
  HS65_LLS_XOR3X2 U18221 ( .A(n7), .B(n4410), .C(n4438), .Z(n4437) );
  HS65_LLS_XNOR2X6 U18222 ( .A(w0[8]), .B(n2814), .Z(n4438) );
  HS65_LL_OAI22X6 U18223 ( .A(n5969), .B(n9130), .C(n9124), .D(n5970), .Z(N210) );
  HS65_LLS_XNOR2X6 U18224 ( .A(w1[24]), .B(text_in_r[88]), .Z(n5969) );
  HS65_LLS_XOR3X2 U18225 ( .A(n5968), .B(n5971), .C(n5972), .Z(n5970) );
  HS65_LLS_XNOR2X6 U18226 ( .A(w1[24]), .B(n529), .Z(n5972) );
  HS65_LL_OAI22X6 U18227 ( .A(n6001), .B(n9129), .C(n9123), .D(n6002), .Z(N194) );
  HS65_LLS_XNOR2X6 U18228 ( .A(w1[16]), .B(text_in_r[80]), .Z(n6001) );
  HS65_LLS_XOR3X2 U18229 ( .A(n5986), .B(n6003), .C(n6004), .Z(n6002) );
  HS65_LLS_XNOR2X6 U18230 ( .A(w1[16]), .B(n50), .Z(n6004) );
  HS65_LL_OAI22X6 U18231 ( .A(n5973), .B(n9130), .C(n9124), .D(n5974), .Z(N201) );
  HS65_LLS_XNOR2X6 U18232 ( .A(w1[23]), .B(text_in_r[87]), .Z(n5973) );
  HS65_LLS_XOR3X2 U18233 ( .A(n52), .B(n5944), .C(n5975), .Z(n5974) );
  HS65_LLS_XNOR2X6 U18234 ( .A(w1[23]), .B(n3208), .Z(n5975) );
  HS65_LL_OAI22X6 U18235 ( .A(n7072), .B(n9129), .C(n9122), .D(n7073), .Z(N164) );
  HS65_LLS_XNOR2X6 U18236 ( .A(w1[2]), .B(text_in_r[66]), .Z(n7072) );
  HS65_LLS_XOR3X2 U18237 ( .A(n5962), .B(n6000), .C(n7074), .Z(n7073) );
  HS65_LLS_XNOR2X6 U18238 ( .A(w1[2]), .B(n3008), .Z(n7074) );
  HS65_LL_OAI22X6 U18239 ( .A(n5949), .B(n9130), .C(n9124), .D(n5950), .Z(N214) );
  HS65_LLS_XNOR2X6 U18240 ( .A(w1[28]), .B(text_in_r[92]), .Z(n5949) );
  HS65_LLS_XOR3X2 U18241 ( .A(n5951), .B(n5952), .C(n5953), .Z(n5950) );
  HS65_LLS_XOR3X2 U18242 ( .A(w1[28]), .B(n2762), .C(n2809), .Z(n5953) );
  HS65_LL_OAI22X6 U18243 ( .A(n5984), .B(n9130), .C(n9124), .D(n5985), .Z(N198) );
  HS65_LLS_XNOR2X6 U18244 ( .A(w1[20]), .B(text_in_r[84]), .Z(n5984) );
  HS65_LLS_XOR3X2 U18245 ( .A(n5986), .B(n5987), .C(n5988), .Z(n5985) );
  HS65_LLS_XOR3X2 U18246 ( .A(w1[20]), .B(n5957), .C(n2786), .Z(n5987) );
  HS65_LL_OAI22X6 U18247 ( .A(n5993), .B(n9130), .C(n9124), .D(n5994), .Z(N196) );
  HS65_LLS_XNOR2X6 U18248 ( .A(w1[18]), .B(text_in_r[82]), .Z(n5993) );
  HS65_LLS_XOR3X2 U18249 ( .A(n5965), .B(n5995), .C(n5996), .Z(n5994) );
  HS65_LLS_XNOR2X6 U18250 ( .A(w1[18]), .B(n2784), .Z(n5996) );
  HS65_LL_OAI22X6 U18251 ( .A(n7597), .B(n9132), .C(n9125), .D(n7598), .Z(N120) );
  HS65_LLS_XNOR2X6 U18252 ( .A(w2[14]), .B(text_in_r[46]), .Z(n7597) );
  HS65_LLS_XOR3X2 U18253 ( .A(n2804), .B(n7568), .C(n7599), .Z(n7598) );
  HS65_LLS_XOR3X2 U18254 ( .A(n2755), .B(w2[14]), .C(n2779), .Z(n7599) );
  HS65_LL_OAI22X6 U18255 ( .A(n6025), .B(n9129), .C(n9123), .D(n6026), .Z(N179) );
  HS65_LLS_XNOR2X6 U18256 ( .A(w1[9]), .B(text_in_r[73]), .Z(n6025) );
  HS65_LLS_XOR3X2 U18257 ( .A(n6000), .B(n6027), .C(n6028), .Z(n6026) );
  HS65_LLS_XNOR2X6 U18258 ( .A(n2807), .B(n52), .Z(n6027) );
  HS65_LL_OAI22X6 U18259 ( .A(n7153), .B(n9129), .C(n9122), .D(n7154), .Z(N163) );
  HS65_LLS_XNOR2X6 U18260 ( .A(w1[1]), .B(text_in_r[65]), .Z(n7153) );
  HS65_LLS_XOR3X2 U18261 ( .A(n6003), .B(n7155), .C(n6396), .Z(n7154) );
  HS65_LLS_XNOR3X2 U18262 ( .A(w1[1]), .B(n5965), .C(n3007), .Z(n7155) );
  HS65_LL_OAI22X6 U18263 ( .A(n8474), .B(n9133), .C(n9128), .D(n8475), .Z(N101) );
  HS65_LLS_XNOR2X6 U18264 ( .A(w2[3]), .B(text_in_r[35]), .Z(n8474) );
  HS65_LLS_XOR3X2 U18265 ( .A(n7550), .B(n8476), .C(n7585), .Z(n8475) );
  HS65_LLS_XNOR3X2 U18266 ( .A(w2[3]), .B(n2616), .C(n3001), .Z(n8476) );
  HS65_LL_OAI22X6 U18267 ( .A(n7556), .B(n9131), .C(n9124), .D(n7557), .Z(N147) );
  HS65_LLS_XNOR2X6 U18268 ( .A(w2[25]), .B(text_in_r[57]), .Z(n7556) );
  HS65_LLS_XOR2X6 U18269 ( .A(n7558), .B(n7559), .Z(n7557) );
  HS65_LLS_XOR3X2 U18270 ( .A(w2[25]), .B(n2898), .C(n2798), .Z(n7558) );
  HS65_LL_OAI22X6 U18271 ( .A(n4421), .B(n9135), .C(n9125), .D(n4422), .Z(N246) );
  HS65_LLS_XNOR2X6 U18272 ( .A(w0[12]), .B(text_in_r[108]), .Z(n4421) );
  HS65_LLS_XOR3X2 U18273 ( .A(n4423), .B(n4395), .C(n4424), .Z(n4422) );
  HS65_LLS_XOR3X2 U18274 ( .A(w0[12]), .B(n2769), .C(n2793), .Z(n4424) );
  HS65_LL_OAI22X6 U18275 ( .A(n2621), .B(n9132), .C(n9124), .D(n2622), .Z(N98)
         );
  HS65_LLS_XNOR2X6 U18276 ( .A(w2[0]), .B(text_in_r[32]), .Z(n2621) );
  HS65_LLS_XOR3X2 U18277 ( .A(n2616), .B(n2623), .C(n2624), .Z(n2622) );
  HS65_LLS_XNOR2X6 U18278 ( .A(w2[0]), .B(n315), .Z(n2624) );
  HS65_LL_OAI22X6 U18279 ( .A(n7929), .B(n9132), .C(n9124), .D(n7930), .Z(N104) );
  HS65_LLS_XNOR2X6 U18280 ( .A(w2[6]), .B(text_in_r[38]), .Z(n7929) );
  HS65_LLS_XOR3X2 U18281 ( .A(n7535), .B(n7572), .C(n7931), .Z(n7930) );
  HS65_LLS_XNOR2X6 U18282 ( .A(w2[6]), .B(n3004), .Z(n7931) );
  HS65_LL_OAI22X6 U18283 ( .A(n6029), .B(n9129), .C(n9123), .D(n6030), .Z(N178) );
  HS65_LLS_XNOR2X6 U18284 ( .A(w1[8]), .B(text_in_r[72]), .Z(n6029) );
  HS65_LLS_XOR3X2 U18285 ( .A(n52), .B(n6003), .C(n6031), .Z(n6030) );
  HS65_LLS_XNOR2X6 U18286 ( .A(w1[8]), .B(n2806), .Z(n6031) );
  HS65_LL_OAI22X6 U18287 ( .A(n4380), .B(n9133), .C(n9126), .D(n4381), .Z(N265) );
  HS65_LLS_XNOR2X6 U18288 ( .A(w0[23]), .B(text_in_r[119]), .Z(n4380) );
  HS65_LLS_XOR3X2 U18289 ( .A(n7), .B(n4351), .C(n4382), .Z(n4381) );
  HS65_LLS_XNOR2X6 U18290 ( .A(w0[23]), .B(n3533), .Z(n4382) );
  HS65_LL_OAI22X6 U18291 ( .A(n7775), .B(n9132), .C(n9123), .D(n7776), .Z(N105) );
  HS65_LLS_XNOR2X6 U18292 ( .A(w2[7]), .B(text_in_r[39]), .Z(n7775) );
  HS65_LLS_XOR3X2 U18293 ( .A(n7546), .B(n7568), .C(n7777), .Z(n7776) );
  HS65_LLS_XNOR2X6 U18294 ( .A(w2[7]), .B(n2781), .Z(n7777) );
  HS65_LL_OAI22X6 U18295 ( .A(n7583), .B(n9133), .C(n9123), .D(n7584), .Z(N132) );
  HS65_LLS_XNOR2X6 U18296 ( .A(w2[18]), .B(text_in_r[50]), .Z(n7583) );
  HS65_LLS_XOR3X2 U18297 ( .A(n2618), .B(n7585), .C(n7586), .Z(n7584) );
  HS65_LLS_XNOR2X6 U18298 ( .A(w2[18]), .B(n2776), .Z(n7586) );
  HS65_LL_OAI22X6 U18299 ( .A(n4356), .B(n9135), .C(n9126), .D(n4357), .Z(N278) );
  HS65_LLS_XNOR2X6 U18300 ( .A(w0[28]), .B(text_in_r[124]), .Z(n4356) );
  HS65_LLS_XOR3X2 U18301 ( .A(n4358), .B(n4359), .C(n4360), .Z(n4357) );
  HS65_LLS_XOR3X2 U18302 ( .A(w0[28]), .B(n2770), .C(n2817), .Z(n4360) );
  HS65_LL_OAI22X6 U18303 ( .A(n4391), .B(n9134), .C(n9126), .D(n4392), .Z(N262) );
  HS65_LLS_XNOR2X6 U18304 ( .A(w0[20]), .B(text_in_r[116]), .Z(n4391) );
  HS65_LLS_XOR3X2 U18305 ( .A(n4393), .B(n4394), .C(n4395), .Z(n4392) );
  HS65_LLS_XOR3X2 U18306 ( .A(w0[20]), .B(n4364), .C(n2794), .Z(n4394) );
  HS65_LL_OAI22X6 U18307 ( .A(n4376), .B(n9135), .C(n9126), .D(n4377), .Z(N274) );
  HS65_LLS_XNOR2X6 U18308 ( .A(w0[24]), .B(text_in_r[120]), .Z(n4376) );
  HS65_LLS_XOR3X2 U18309 ( .A(n4375), .B(n4378), .C(n4379), .Z(n4377) );
  HS65_LLS_XNOR2X6 U18310 ( .A(w0[24]), .B(n2766), .Z(n4379) );
  HS65_LL_OAI22X6 U18311 ( .A(n4408), .B(n9133), .C(n9125), .D(n4409), .Z(N258) );
  HS65_LLS_XNOR2X6 U18312 ( .A(w0[16]), .B(text_in_r[112]), .Z(n4408) );
  HS65_LLS_XOR3X2 U18313 ( .A(n4393), .B(n4410), .C(n4411), .Z(n4409) );
  HS65_LLS_XNOR2X6 U18314 ( .A(w0[16]), .B(n2790), .Z(n4411) );
  HS65_LL_OAI22X6 U18315 ( .A(n4400), .B(n9135), .C(n9122), .D(n4401), .Z(N260) );
  HS65_LLS_XNOR2X6 U18316 ( .A(w0[18]), .B(text_in_r[114]), .Z(n4400) );
  HS65_LLS_XOR3X2 U18317 ( .A(n4372), .B(n4402), .C(n4403), .Z(n4401) );
  HS65_LLS_XNOR2X6 U18318 ( .A(w0[18]), .B(n2792), .Z(n4403) );
  HS65_LL_AND2X4 U18319 ( .A(sa03[0]), .B(sa03[1]), .Z(n4147) );
  HS65_LL_AND2X4 U18320 ( .A(sa02[2]), .B(n357), .Z(n8931) );
  HS65_LL_AND2X4 U18321 ( .A(sa31[2]), .B(n401), .Z(n8986) );
  HS65_LL_AND2X4 U18322 ( .A(sa13[1]), .B(sa13[0]), .Z(n9106) );
  HS65_LL_AND2X4 U18323 ( .A(sa20[1]), .B(sa20[0]), .Z(n9048) );
  HS65_LL_OAI22X6 U18324 ( .A(n4429), .B(n9133), .C(n9126), .D(n4430), .Z(N244) );
  HS65_LLS_XNOR2X6 U18325 ( .A(w0[10]), .B(text_in_r[106]), .Z(n4429) );
  HS65_LLS_XNOR3X2 U18326 ( .A(n2816), .B(n4431), .C(n4402), .Z(n4430) );
  HS65_LLS_XOR3X2 U18327 ( .A(n2767), .B(n947), .C(n229), .Z(n4431) );
  HS65_LLS_XOR3X2 U18328 ( .A(n1374), .B(\u0/rcon [26]), .C(n958), .Z(n982) );
  HS65_LL_NOR4ABX2 U18329 ( .A(n1375), .B(n1376), .C(n1377), .D(n1378), .Z(
        n1374) );
  HS65_LL_CBI4I1X5 U18330 ( .A(n1163), .B(n1111), .C(n1145), .D(n1341), .Z(
        n1378) );
  HS65_LL_AOI212X4 U18331 ( .A(n852), .B(n871), .C(n860), .D(n1123), .E(n1393), 
        .Z(n1376) );
  HS65_LLS_XOR3X2 U18332 ( .A(n957), .B(\u0/rcon [25]), .C(n1396), .Z(n983) );
  HS65_LL_NAND4ABX3 U18333 ( .A(n1397), .B(n1398), .C(n1399), .D(n1400), .Z(
        n1396) );
  HS65_LL_CB4I6X9 U18334 ( .A(n844), .B(n849), .C(n871), .D(n1334), .Z(n1397)
         );
  HS65_LL_AOI222X2 U18335 ( .A(n863), .B(n841), .C(n860), .D(n1419), .E(n872), 
        .F(n840), .Z(n1399) );
  HS65_LLS_XOR3X2 U18336 ( .A(n961), .B(\u0/rcon [30]), .C(n1132), .Z(n978) );
  HS65_LL_NAND4ABX3 U18337 ( .A(n1133), .B(n1134), .C(n1135), .D(n1136), .Z(
        n1132) );
  HS65_LL_AOI212X4 U18338 ( .A(n873), .B(n839), .C(n870), .D(n851), .E(n1142), 
        .Z(n1135) );
  HS65_LL_CBI4I1X5 U18339 ( .A(n1148), .B(n1110), .C(n1149), .D(n1150), .Z(
        n1133) );
  HS65_LL_IVX9 U18340 ( .A(sa22[4]), .Z(n249) );
  HS65_LL_IVX9 U18341 ( .A(sa11[4]), .Z(n466) );
  HS65_LL_IVX9 U18342 ( .A(sa33[6]), .Z(n26) );
  HS65_LL_IVX9 U18343 ( .A(sa33[4]), .Z(n27) );
  HS65_LL_IVX9 U18344 ( .A(sa00[4]), .Z(n682) );
  HS65_LL_IVX9 U18345 ( .A(sa12[4]), .Z(n291) );
  HS65_LL_IVX9 U18346 ( .A(sa01[4]), .Z(n506) );
  HS65_LL_IVX9 U18347 ( .A(sa30[6]), .Z(n548) );
  HS65_LL_IVX9 U18348 ( .A(sa30[4]), .Z(n549) );
  HS65_LL_IVX9 U18349 ( .A(sa23[6]), .Z(n70) );
  HS65_LL_IVX9 U18350 ( .A(sa23[4]), .Z(n71) );
  HS65_LL_IVX9 U18351 ( .A(sa11[6]), .Z(n465) );
  HS65_LL_IVX9 U18352 ( .A(sa00[6]), .Z(n681) );
  HS65_LL_IVX9 U18353 ( .A(sa22[6]), .Z(n248) );
  HS65_LL_IVX9 U18354 ( .A(sa12[6]), .Z(n290) );
  HS65_LL_IVX9 U18355 ( .A(sa01[6]), .Z(n505) );
  HS65_LL_IVX9 U18356 ( .A(sa22[0]), .Z(n271) );
  HS65_LL_IVX9 U18357 ( .A(sa11[0]), .Z(n488) );
  HS65_LL_IVX9 U18358 ( .A(sa33[0]), .Z(n49) );
  HS65_LL_IVX9 U18359 ( .A(sa00[0]), .Z(n704) );
  HS65_LL_IVX9 U18360 ( .A(sa12[0]), .Z(n313) );
  HS65_LL_IVX9 U18361 ( .A(sa01[0]), .Z(n528) );
  HS65_LL_IVX9 U18362 ( .A(sa30[0]), .Z(n571) );
  HS65_LL_IVX9 U18363 ( .A(sa23[0]), .Z(n93) );
  HS65_LL_IVX9 U18364 ( .A(sa20[0]), .Z(n619) );
  HS65_LL_IVX9 U18365 ( .A(sa13[0]), .Z(n139) );
  HS65_LL_OAI22X6 U18366 ( .A(n756), .B(n9145), .C(n1072), .D(n9137), .Z(
        \u0/N174 ) );
  HS65_LL_IVX9 U18367 ( .A(key[32]), .Z(n756) );
  HS65_LL_OAI22X6 U18368 ( .A(n748), .B(n9145), .C(n1056), .D(n9138), .Z(
        \u0/N182 ) );
  HS65_LL_IVX9 U18369 ( .A(key[40]), .Z(n748) );
  HS65_LL_OAI22X6 U18370 ( .A(n753), .B(n9145), .C(n1066), .D(n9137), .Z(
        \u0/N177 ) );
  HS65_LL_IVX9 U18371 ( .A(key[35]), .Z(n753) );
  HS65_LL_OAI22X6 U18372 ( .A(n744), .B(n9145), .C(n1048), .D(n9138), .Z(
        \u0/N186 ) );
  HS65_LL_IVX9 U18373 ( .A(key[44]), .Z(n744) );
  HS65_LL_OAI22X6 U18374 ( .A(n728), .B(n9145), .C(n1016), .D(n9139), .Z(
        \u0/N202 ) );
  HS65_LL_IVX9 U18375 ( .A(key[60]), .Z(n728) );
  HS65_LL_OAI22X6 U18376 ( .A(n740), .B(n9148), .C(n1040), .D(n9139), .Z(
        \u0/N190 ) );
  HS65_LL_IVX9 U18377 ( .A(key[48]), .Z(n740) );
  HS65_LL_OAI22X6 U18378 ( .A(n732), .B(n9148), .C(n1024), .D(n9139), .Z(
        \u0/N198 ) );
  HS65_LL_IVX9 U18379 ( .A(key[56]), .Z(n732) );
  HS65_LL_OAI22X6 U18380 ( .A(n746), .B(n9149), .C(n1052), .D(n9138), .Z(
        \u0/N184 ) );
  HS65_LL_IVX9 U18381 ( .A(key[42]), .Z(n746) );
  HS65_LL_OAI22X6 U18382 ( .A(n749), .B(n9148), .C(n1058), .D(n9138), .Z(
        \u0/N181 ) );
  HS65_LL_IVX9 U18383 ( .A(key[39]), .Z(n749) );
  HS65_LL_OAI22X6 U18384 ( .A(n747), .B(n9143), .C(n1054), .D(n9138), .Z(
        \u0/N183 ) );
  HS65_LL_IVX9 U18385 ( .A(key[41]), .Z(n747) );
  HS65_LL_OAI22X6 U18386 ( .A(n754), .B(n9149), .C(n1068), .D(n9137), .Z(
        \u0/N176 ) );
  HS65_LL_IVX9 U18387 ( .A(key[34]), .Z(n754) );
  HS65_LL_OAI22X6 U18388 ( .A(n741), .B(n9148), .C(n1042), .D(n9139), .Z(
        \u0/N189 ) );
  HS65_LL_IVX9 U18389 ( .A(key[47]), .Z(n741) );
  HS65_LL_OAI22X6 U18390 ( .A(n739), .B(n9148), .C(n1038), .D(n9139), .Z(
        \u0/N191 ) );
  HS65_LL_IVX9 U18391 ( .A(key[49]), .Z(n739) );
  HS65_LL_OAI22X6 U18392 ( .A(n750), .B(n9118), .C(n1060), .D(n9137), .Z(
        \u0/N180 ) );
  HS65_LL_IVX9 U18393 ( .A(key[38]), .Z(n750) );
  HS65_LL_OAI22X6 U18394 ( .A(n745), .B(n9143), .C(n1050), .D(n9138), .Z(
        \u0/N185 ) );
  HS65_LL_IVX9 U18395 ( .A(key[43]), .Z(n745) );
  HS65_LL_OAI22X6 U18396 ( .A(n726), .B(n9148), .C(n1012), .D(n9139), .Z(
        \u0/N204 ) );
  HS65_LL_IVX9 U18397 ( .A(key[62]), .Z(n726) );
  HS65_LL_OAI22X6 U18398 ( .A(n752), .B(n9118), .C(n1064), .D(n9137), .Z(
        \u0/N178 ) );
  HS65_LL_IVX9 U18399 ( .A(key[36]), .Z(n752) );
  HS65_LL_OAI22X6 U18400 ( .A(n743), .B(n9148), .C(n1046), .D(n9138), .Z(
        \u0/N187 ) );
  HS65_LL_IVX9 U18401 ( .A(key[45]), .Z(n743) );
  HS65_LL_OAI22X6 U18402 ( .A(n735), .B(n9148), .C(n1030), .D(n9139), .Z(
        \u0/N195 ) );
  HS65_LL_IVX9 U18403 ( .A(key[53]), .Z(n735) );
  HS65_LL_OAI22X6 U18404 ( .A(n751), .B(n9118), .C(n1062), .D(n9137), .Z(
        \u0/N179 ) );
  HS65_LL_IVX9 U18405 ( .A(key[37]), .Z(n751) );
  HS65_LL_OAI22X6 U18406 ( .A(n755), .B(n9118), .C(n1070), .D(n9137), .Z(
        \u0/N175 ) );
  HS65_LL_IVX9 U18407 ( .A(key[33]), .Z(n755) );
  HS65_LL_OAI22X6 U18408 ( .A(n742), .B(n9148), .C(n1044), .D(n9139), .Z(
        \u0/N188 ) );
  HS65_LL_IVX9 U18409 ( .A(key[46]), .Z(n742) );
  HS65_LL_OAI22X6 U18410 ( .A(n736), .B(n9144), .C(n1032), .D(n9139), .Z(
        \u0/N194 ) );
  HS65_LL_IVX9 U18411 ( .A(key[52]), .Z(n736) );
  HS65_LL_IVX9 U18412 ( .A(sa10[1]), .Z(n664) );
  HS65_LL_IVX9 U18413 ( .A(sa32[3]), .Z(n222) );
  HS65_LL_IVX9 U18414 ( .A(sa21[3]), .Z(n444) );
  HS65_LL_IVX9 U18415 ( .A(sa31[3]), .Z(n401) );
  HS65_LL_IVX9 U18416 ( .A(sa02[3]), .Z(n357) );
  HS65_LL_IVX9 U18417 ( .A(sa03[1]), .Z(n182) );
  HS65_LL_OAI22X6 U18418 ( .A(n725), .B(n9143), .C(n1010), .D(n9139), .Z(
        \u0/N205 ) );
  HS65_LL_IVX9 U18419 ( .A(key[63]), .Z(n725) );
  HS65_LL_OAI22X6 U18420 ( .A(n733), .B(n9143), .C(n1026), .D(n9139), .Z(
        \u0/N197 ) );
  HS65_LL_IVX9 U18421 ( .A(key[55]), .Z(n733) );
  HS65_LL_OAI22X6 U18422 ( .A(n731), .B(n9143), .C(n1022), .D(n9138), .Z(
        \u0/N199 ) );
  HS65_LL_IVX9 U18423 ( .A(key[57]), .Z(n731) );
  HS65_LL_OAI22X6 U18424 ( .A(n738), .B(n9143), .C(n1036), .D(n9139), .Z(
        \u0/N192 ) );
  HS65_LL_IVX9 U18425 ( .A(key[50]), .Z(n738) );
  HS65_LL_OAI22X6 U18426 ( .A(n729), .B(n9143), .C(n1018), .D(n9138), .Z(
        \u0/N201 ) );
  HS65_LL_IVX9 U18427 ( .A(key[59]), .Z(n729) );
  HS65_LL_OAI22X6 U18428 ( .A(n730), .B(n9143), .C(n1020), .D(n9138), .Z(
        \u0/N200 ) );
  HS65_LL_IVX9 U18429 ( .A(key[58]), .Z(n730) );
  HS65_LL_OAI22X6 U18430 ( .A(n737), .B(n9143), .C(n1034), .D(n9139), .Z(
        \u0/N193 ) );
  HS65_LL_IVX9 U18431 ( .A(key[51]), .Z(n737) );
  HS65_LL_OAI22X6 U18432 ( .A(n727), .B(n9143), .C(n1014), .D(n9138), .Z(
        \u0/N203 ) );
  HS65_LL_IVX9 U18433 ( .A(key[61]), .Z(n727) );
  HS65_LL_OAI22X6 U18434 ( .A(n734), .B(n9143), .C(n1028), .D(n9139), .Z(
        \u0/N196 ) );
  HS65_LL_IVX9 U18435 ( .A(key[54]), .Z(n734) );
  HS65_LLS_XOR3X2 U18436 ( .A(n1105), .B(\u0/rcon [31]), .C(n962), .Z(n977) );
  HS65_LL_NOR3X4 U18437 ( .A(n1106), .B(n1107), .C(n1108), .Z(n1105) );
  HS65_LL_OAI212X5 U18438 ( .A(n1109), .B(n1110), .C(n1111), .D(n1112), .E(
        n1113), .Z(n1108) );
  HS65_LL_NAND4ABX3 U18439 ( .A(n1119), .B(n1120), .C(n1121), .D(n1122), .Z(
        n1107) );
  HS65_LLS_XOR3X2 U18440 ( .A(n1193), .B(\u0/rcon [28]), .C(n960), .Z(n980) );
  HS65_LL_NOR3X4 U18441 ( .A(n1194), .B(n1195), .C(n1196), .Z(n1193) );
  HS65_LL_OAI212X5 U18442 ( .A(n1197), .B(n1112), .C(n1198), .D(n1199), .E(
        n1200), .Z(n1196) );
  HS65_LL_NAND4ABX3 U18443 ( .A(n1201), .B(n1202), .C(n1203), .D(n1204), .Z(
        n1195) );
  HS65_LLS_XOR3X2 U18444 ( .A(n956), .B(\u0/rcon [24]), .C(n1421), .Z(n984) );
  HS65_LL_NAND4ABX3 U18445 ( .A(n1422), .B(n1423), .C(n1424), .D(n1425), .Z(
        n1421) );
  HS65_LL_MX41X7 U18446 ( .D0(n852), .S0(n869), .D1(n853), .S1(n861), .D2(n872), .S2(n845), .D3(n873), .S3(n1185), .Z(n1423) );
  HS65_LL_NOR4ABX2 U18447 ( .A(n1183), .B(n1318), .C(n1426), .D(n1332), .Z(
        n1425) );
  HS65_LLS_XOR3X2 U18448 ( .A(n959), .B(\u0/rcon [27]), .C(n1255), .Z(n981) );
  HS65_LL_NAND4ABX3 U18449 ( .A(n1256), .B(n1257), .C(n1258), .D(n1259), .Z(
        n1255) );
  HS65_LL_AOI212X4 U18450 ( .A(n855), .B(n1260), .C(n871), .D(n1237), .E(n1261), .Z(n1259) );
  HS65_LL_MX41X7 U18451 ( .D0(n842), .S0(n866), .D1(n870), .S1(n854), .D2(n840), .S2(n861), .D3(n872), .S3(n1185), .Z(n1257) );
  HS65_LL_AND2X4 U18452 ( .A(sa21[2]), .B(sa21[3]), .Z(n4325) );
  HS65_LL_AND2X4 U18453 ( .A(sa02[2]), .B(sa02[3]), .Z(n8916) );
  HS65_LL_AND2X4 U18454 ( .A(sa20[1]), .B(n619), .Z(n9045) );
  HS65_LL_AND2X4 U18455 ( .A(sa13[1]), .B(n139), .Z(n9103) );
  HS65_LL_AND2X4 U18456 ( .A(sa11[1]), .B(n488), .Z(n5920) );
  HS65_LL_AND2X4 U18457 ( .A(sa22[1]), .B(n271), .Z(n5861) );
  HS65_LL_AND2X4 U18458 ( .A(sa12[1]), .B(n313), .Z(n7512) );
  HS65_LL_AND2X4 U18459 ( .A(sa33[1]), .B(n49), .Z(n5750) );
  HS65_LL_AND2X4 U18460 ( .A(sa00[1]), .B(n704), .Z(n5812) );
  HS65_LL_AND2X4 U18461 ( .A(sa01[1]), .B(n528), .Z(n7404) );
  HS65_LL_AND2X4 U18462 ( .A(sa30[1]), .B(n571), .Z(n7342) );
  HS65_LL_AND2X4 U18463 ( .A(sa23[1]), .B(n93), .Z(n7454) );
  HS65_LL_AND2X4 U18464 ( .A(sa21[2]), .B(n444), .Z(n4339) );
  HS65_LL_AND2X4 U18465 ( .A(sa32[2]), .B(n222), .Z(n4210) );
  HS65_LL_AND2X4 U18466 ( .A(sa33[1]), .B(sa33[0]), .Z(n5728) );
  HS65_LL_AND2X4 U18467 ( .A(sa30[1]), .B(sa30[0]), .Z(n7320) );
  HS65_LL_AND2X4 U18468 ( .A(sa10[0]), .B(n664), .Z(n4281) );
  HS65_LL_AND2X4 U18469 ( .A(sa03[0]), .B(n182), .Z(n4155) );
  HS65_LLS_XNOR2X6 U18470 ( .A(w0[6]), .B(n2260), .Z(n1002) );
  HS65_LL_NAND4ABX3 U18471 ( .A(n2261), .B(n2262), .C(n2263), .D(n2264), .Z(
        n2260) );
  HS65_LL_AOI212X4 U18472 ( .A(n914), .B(n880), .C(n911), .D(n892), .E(n2270), 
        .Z(n2263) );
  HS65_LL_CBI4I1X5 U18473 ( .A(n2272), .B(n2273), .C(n2274), .D(n2275), .Z(
        n2262) );
  HS65_LL_OAI22X6 U18474 ( .A(n2719), .B(n9131), .C(n9128), .D(n2720), .Z(N57)
         );
  HS65_LLS_XNOR2X6 U18475 ( .A(w3[15]), .B(text_in_r[15]), .Z(n2719) );
  HS65_LLS_XOR3X2 U18476 ( .A(n2637), .B(n2654), .C(n2721), .Z(n2720) );
  HS65_LLS_XOR3X2 U18477 ( .A(n2722), .B(w3[15]), .C(n2687), .Z(n2721) );
  HS65_LLS_XOR3X2 U18478 ( .A(n574), .B(w2[10]), .C(n2751), .Z(n7613) );
  HS65_LL_OAI22X6 U18479 ( .A(n2625), .B(n9132), .C(n9128), .D(n2626), .Z(N89)
         );
  HS65_LLS_XNOR2X6 U18480 ( .A(w3[31]), .B(text_in_r[31]), .Z(n2625) );
  HS65_LLS_XOR3X2 U18481 ( .A(n2627), .B(n2628), .C(n2629), .Z(n2626) );
  HS65_LLS_XOR3X2 U18482 ( .A(n2630), .B(w3[31]), .C(n2631), .Z(n2629) );
  HS65_LL_OAI22X6 U18483 ( .A(n7529), .B(n9129), .C(n9122), .D(n7530), .Z(N153) );
  HS65_LLS_XNOR2X6 U18484 ( .A(w2[31]), .B(text_in_r[63]), .Z(n7529) );
  HS65_LLS_XNOR3X2 U18485 ( .A(n3004), .B(n7531), .C(n7532), .Z(n7530) );
  HS65_LLS_XOR3X2 U18486 ( .A(n2804), .B(w2[31]), .C(n2805), .Z(n7531) );
  HS65_LL_OAI22X6 U18487 ( .A(n7701), .B(n9132), .C(n9122), .D(n7702), .Z(N114) );
  HS65_LLS_XNOR2X6 U18488 ( .A(w2[8]), .B(text_in_r[40]), .Z(n7701) );
  HS65_LLS_XOR3X2 U18489 ( .A(n2619), .B(n7532), .C(n7703), .Z(n7702) );
  HS65_LLS_XNOR2X6 U18490 ( .A(w2[8]), .B(n2798), .Z(n7703) );
  HS65_LLS_XOR3X2 U18491 ( .A(n2758), .B(w1[9]), .C(n2782), .Z(n6028) );
  HS65_LL_AND2X4 U18492 ( .A(sa32[2]), .B(sa32[3]), .Z(n4216) );
  HS65_LL_AND2X4 U18493 ( .A(sa31[2]), .B(sa31[3]), .Z(n8984) );
  HS65_LL_OAI22X6 U18494 ( .A(n2679), .B(n9131), .C(n9128), .D(n2680), .Z(N73)
         );
  HS65_LLS_XNOR2X6 U18495 ( .A(w3[23]), .B(text_in_r[23]), .Z(n2679) );
  HS65_LLS_XOR3X2 U18496 ( .A(n2628), .B(n2636), .C(n2681), .Z(n2680) );
  HS65_LLS_XNOR2X6 U18497 ( .A(w3[23]), .B(n2682), .Z(n2681) );
  HS65_LL_OAI22X6 U18498 ( .A(n2746), .B(n9136), .C(n9127), .D(n2747), .Z(N50)
         );
  HS65_LLS_XNOR2X6 U18499 ( .A(w3[8]), .B(text_in_r[8]), .Z(n2746) );
  HS65_LLS_XOR3X2 U18500 ( .A(n2628), .B(n2716), .C(n2748), .Z(n2747) );
  HS65_LLS_XNOR2X6 U18501 ( .A(w3[8]), .B(n2672), .Z(n2748) );
  HS65_LL_OAI22X6 U18502 ( .A(n7591), .B(n9129), .C(n9122), .D(n7592), .Z(N130) );
  HS65_LLS_XNOR2X6 U18503 ( .A(w2[16]), .B(text_in_r[48]), .Z(n7591) );
  HS65_LLS_XOR3X2 U18504 ( .A(n2619), .B(n7576), .C(n7593), .Z(n7592) );
  HS65_LLS_XNOR2X6 U18505 ( .A(w2[16]), .B(n2774), .Z(n7593) );
  HS65_LL_OAI22X6 U18506 ( .A(n4396), .B(n9135), .C(n9125), .D(n4397), .Z(N261) );
  HS65_LLS_XNOR2X6 U18507 ( .A(w0[19]), .B(text_in_r[115]), .Z(n4396) );
  HS65_LLS_XOR3X2 U18508 ( .A(n4393), .B(n4398), .C(n4399), .Z(n4397) );
  HS65_LLS_XOR3X2 U18509 ( .A(w0[19]), .B(n4369), .C(n2793), .Z(n4398) );
  HS65_LL_OAI22X6 U18510 ( .A(n6008), .B(n9129), .C(n9123), .D(n6009), .Z(N184) );
  HS65_LLS_XNOR2X6 U18511 ( .A(w1[14]), .B(text_in_r[78]), .Z(n6008) );
  HS65_LLS_XOR3X2 U18512 ( .A(n2812), .B(n5978), .C(n6010), .Z(n6009) );
  HS65_LLS_XOR3X2 U18513 ( .A(n2763), .B(w1[14]), .C(n2787), .Z(n6010) );
  HS65_LL_OAI22X6 U18514 ( .A(n4415), .B(n9135), .C(n9122), .D(n4416), .Z(N248) );
  HS65_LLS_XNOR2X6 U18515 ( .A(w0[14]), .B(text_in_r[110]), .Z(n4415) );
  HS65_LLS_XOR3X2 U18516 ( .A(n2820), .B(n4385), .C(n4417), .Z(n4416) );
  HS65_LLS_XOR3X2 U18517 ( .A(n2771), .B(n948), .C(n2795), .Z(n4417) );
  HS65_LL_OAI22X6 U18518 ( .A(n5976), .B(n9130), .C(n9124), .D(n5977), .Z(N200) );
  HS65_LLS_XNOR2X6 U18519 ( .A(w1[22]), .B(text_in_r[86]), .Z(n5976) );
  HS65_LLS_XOR3X2 U18520 ( .A(n5948), .B(n5978), .C(n5979), .Z(n5977) );
  HS65_LLS_XNOR2X6 U18521 ( .A(w1[22]), .B(n53), .Z(n5979) );
  HS65_LL_OAI22X6 U18522 ( .A(n4383), .B(n9133), .C(n9126), .D(n4384), .Z(N264) );
  HS65_LLS_XNOR2X6 U18523 ( .A(w0[22]), .B(text_in_r[118]), .Z(n4383) );
  HS65_LLS_XOR3X2 U18524 ( .A(n4355), .B(n4385), .C(n4386), .Z(n4384) );
  HS65_LLS_XNOR2X6 U18525 ( .A(w0[22]), .B(n231), .Z(n4386) );
  HS65_LL_OAI22X6 U18526 ( .A(n6032), .B(n9129), .C(n9123), .D(n6033), .Z(N169) );
  HS65_LLS_XNOR2X6 U18527 ( .A(w1[7]), .B(text_in_r[71]), .Z(n6032) );
  HS65_LLS_XOR3X2 U18528 ( .A(n5968), .B(n5978), .C(n6034), .Z(n6033) );
  HS65_LLS_XNOR2X6 U18529 ( .A(w1[7]), .B(n2789), .Z(n6034) );
  HS65_LL_OAI22X6 U18530 ( .A(n4439), .B(n9133), .C(n9125), .D(n4440), .Z(N233) );
  HS65_LLS_XNOR2X6 U18531 ( .A(w0[7]), .B(text_in_r[103]), .Z(n4439) );
  HS65_LLS_XOR3X2 U18532 ( .A(n4375), .B(n4385), .C(n4441), .Z(n4440) );
  HS65_LLS_XNOR2X6 U18533 ( .A(w0[7]), .B(n2797), .Z(n4441) );
  HS65_LL_OAI22X6 U18534 ( .A(n4412), .B(n9134), .C(n9126), .D(n4413), .Z(N249) );
  HS65_LLS_XNOR2X6 U18535 ( .A(w0[15]), .B(text_in_r[111]), .Z(n4412) );
  HS65_LLS_XOR3X2 U18536 ( .A(n2796), .B(n4414), .C(n4375), .Z(n4413) );
  HS65_LLS_XOR3X2 U18537 ( .A(n2772), .B(n949), .C(n2773), .Z(n4414) );
  HS65_LL_OAI22X6 U18538 ( .A(n6005), .B(n9129), .C(n9123), .D(n6006), .Z(N185) );
  HS65_LLS_XNOR2X6 U18539 ( .A(w1[15]), .B(text_in_r[79]), .Z(n6005) );
  HS65_LLS_XOR3X2 U18540 ( .A(n2788), .B(n6007), .C(n5968), .Z(n6006) );
  HS65_LLS_XOR3X2 U18541 ( .A(n2764), .B(n934), .C(n2765), .Z(n6007) );
  HS65_LL_OAI22X6 U18542 ( .A(n7587), .B(n9136), .C(n9127), .D(n7588), .Z(N131) );
  HS65_LLS_XNOR2X6 U18543 ( .A(w2[17]), .B(text_in_r[49]), .Z(n7587) );
  HS65_LLS_XOR3X2 U18544 ( .A(n7576), .B(n7589), .C(n7590), .Z(n7588) );
  HS65_LLS_XOR3X2 U18545 ( .A(w2[17]), .B(n2623), .C(n2775), .Z(n7589) );
  HS65_LL_OAI22X6 U18546 ( .A(n4361), .B(n9134), .C(n9126), .D(n4362), .Z(N277) );
  HS65_LLS_XNOR2X6 U18547 ( .A(w0[27]), .B(text_in_r[123]), .Z(n4361) );
  HS65_LLS_XOR3X2 U18548 ( .A(n4363), .B(n4364), .C(n4365), .Z(n4362) );
  HS65_LLS_XOR3X2 U18549 ( .A(n959), .B(n2769), .C(n2816), .Z(n4365) );
  HS65_LL_OAI22X6 U18550 ( .A(n2723), .B(n9131), .C(n9128), .D(n2724), .Z(N56)
         );
  HS65_LLS_XNOR2X6 U18551 ( .A(w3[14]), .B(text_in_r[14]), .Z(n2723) );
  HS65_LLS_XOR3X2 U18552 ( .A(n2644), .B(n2725), .C(n2685), .Z(n2724) );
  HS65_LLS_XOR3X2 U18553 ( .A(n2627), .B(n837), .C(n2692), .Z(n2725) );
  HS65_LL_OAI22X6 U18554 ( .A(n2632), .B(n9132), .C(n9127), .D(n2633), .Z(N88)
         );
  HS65_LLS_XNOR2X6 U18555 ( .A(w3[30]), .B(text_in_r[30]), .Z(n2632) );
  HS65_LLS_XOR3X2 U18556 ( .A(n2634), .B(n2635), .C(n2636), .Z(n2633) );
  HS65_LLS_XOR3X2 U18557 ( .A(n2637), .B(n919), .C(n2638), .Z(n2635) );
  HS65_LL_OAI22X6 U18558 ( .A(n2709), .B(n9131), .C(n9128), .D(n2710), .Z(N67)
         );
  HS65_LLS_XNOR2X6 U18559 ( .A(w3[17]), .B(text_in_r[17]), .Z(n2709) );
  HS65_LLS_XOR3X2 U18560 ( .A(n2695), .B(n2711), .C(n2712), .Z(n2710) );
  HS65_LLS_XOR3X2 U18561 ( .A(n857), .B(n2677), .C(n2713), .Z(n2711) );
  HS65_LL_OAI22X6 U18562 ( .A(n5561), .B(n9130), .C(n9125), .D(n5562), .Z(N227) );
  HS65_LLS_XNOR2X6 U18563 ( .A(w0[1]), .B(text_in_r[97]), .Z(n5561) );
  HS65_LLS_XOR3X2 U18564 ( .A(n4410), .B(n5563), .C(n4803), .Z(n5562) );
  HS65_LLS_XOR3X2 U18565 ( .A(n943), .B(n4372), .C(n3210), .Z(n5563) );
  HS65_LL_OAI22X6 U18566 ( .A(n7638), .B(n9132), .C(n9127), .D(n7639), .Z(N115) );
  HS65_LLS_XNOR2X6 U18567 ( .A(w2[9]), .B(text_in_r[41]), .Z(n7638) );
  HS65_LLS_XOR3X2 U18568 ( .A(n7640), .B(n7590), .C(n7641), .Z(n7639) );
  HS65_LLS_XOR3X2 U18569 ( .A(w2[9]), .B(n2799), .C(n2750), .Z(n7641) );
  HS65_LL_OAI22X6 U18570 ( .A(n8842), .B(n9134), .C(n9128), .D(n8843), .Z(N100) );
  HS65_LLS_XNOR2X6 U18571 ( .A(w2[2]), .B(text_in_r[34]), .Z(n8842) );
  HS65_LLS_XOR3X2 U18572 ( .A(n7555), .B(n7590), .C(n8844), .Z(n8843) );
  HS65_LLS_XNOR2X6 U18573 ( .A(w2[2]), .B(n3000), .Z(n8844) );
  HS65_LL_OAI22X6 U18574 ( .A(n2699), .B(n9131), .C(n9128), .D(n2700), .Z(N69)
         );
  HS65_LLS_XNOR2X6 U18575 ( .A(w3[19]), .B(text_in_r[19]), .Z(n2699) );
  HS65_LLS_XOR3X2 U18576 ( .A(n2695), .B(n2701), .C(n2702), .Z(n2700) );
  HS65_LLS_XOR3X2 U18577 ( .A(n859), .B(n2665), .C(n2703), .Z(n2701) );
  HS65_LL_OAI22X6 U18578 ( .A(n7552), .B(n9136), .C(n9122), .D(n7553), .Z(N148) );
  HS65_LLS_XNOR2X6 U18579 ( .A(w2[26]), .B(text_in_r[58]), .Z(n7552) );
  HS65_LLS_XOR3X2 U18580 ( .A(n2752), .B(n7554), .C(n7555), .Z(n7553) );
  HS65_LLS_XOR3X2 U18581 ( .A(n2620), .B(n928), .C(n2799), .Z(n7554) );
  HS65_LL_OAI22X6 U18582 ( .A(n5115), .B(n9130), .C(n9125), .D(n5116), .Z(N229) );
  HS65_LLS_XNOR2X6 U18583 ( .A(w0[3]), .B(text_in_r[99]), .Z(n5115) );
  HS65_LLS_XOR3X2 U18584 ( .A(n4402), .B(n5117), .C(n4803), .Z(n5116) );
  HS65_LLS_XOR3X2 U18585 ( .A(n944), .B(n4364), .C(n3212), .Z(n5117) );
  HS65_LL_OAI22X6 U18586 ( .A(n4800), .B(n9130), .C(n9125), .D(n4801), .Z(N230) );
  HS65_LLS_XNOR2X6 U18587 ( .A(w0[4]), .B(text_in_r[100]), .Z(n4800) );
  HS65_LLS_XOR3X2 U18588 ( .A(n4399), .B(n4802), .C(n4803), .Z(n4801) );
  HS65_LLS_XOR3X2 U18589 ( .A(n945), .B(n4359), .C(n3213), .Z(n4802) );
  HS65_LL_OAI22X6 U18590 ( .A(n3975), .B(n9135), .C(n9126), .D(n3976), .Z(N35)
         );
  HS65_LLS_XNOR2X6 U18591 ( .A(w3[1]), .B(text_in_r[1]), .Z(n3975) );
  HS65_LLS_XOR3X2 U18592 ( .A(n2716), .B(n3977), .C(n3218), .Z(n3976) );
  HS65_LLS_XOR3X2 U18593 ( .A(w3[1]), .B(n2669), .C(n2896), .Z(n3977) );
  HS65_LL_OAI22X6 U18594 ( .A(n3215), .B(n9136), .C(n9127), .D(n3216), .Z(N38)
         );
  HS65_LLS_XNOR2X6 U18595 ( .A(w3[4]), .B(text_in_r[4]), .Z(n3215) );
  HS65_LLS_XOR3X2 U18596 ( .A(n2702), .B(n3217), .C(n3218), .Z(n3216) );
  HS65_LLS_XOR3X2 U18597 ( .A(n794), .B(n2649), .C(n2645), .Z(n3217) );
  HS65_LL_OAI22X6 U18598 ( .A(n3534), .B(n9136), .C(n9127), .D(n3535), .Z(N37)
         );
  HS65_LLS_XNOR2X6 U18599 ( .A(w3[3]), .B(text_in_r[3]), .Z(n3534) );
  HS65_LLS_XOR3X2 U18600 ( .A(n2706), .B(n3536), .C(n3218), .Z(n3535) );
  HS65_LLS_XOR3X2 U18601 ( .A(n777), .B(n2660), .C(n2652), .Z(n3536) );
  HS65_LL_OAI22X6 U18602 ( .A(n5665), .B(n9130), .C(n9125), .D(n5666), .Z(N226) );
  HS65_LLS_XNOR2X6 U18603 ( .A(w0[0]), .B(text_in_r[96]), .Z(n5665) );
  HS65_LLS_XOR3X2 U18604 ( .A(n4378), .B(n4803), .C(n5667), .Z(n5666) );
  HS65_LLS_XNOR2X6 U18605 ( .A(w0[0]), .B(n3209), .Z(n5667) );
  HS65_LL_OAI22X6 U18606 ( .A(n7257), .B(n9129), .C(n9122), .D(n7258), .Z(N162) );
  HS65_LLS_XNOR2X6 U18607 ( .A(w1[0]), .B(text_in_r[64]), .Z(n7257) );
  HS65_LLS_XOR3X2 U18608 ( .A(n5971), .B(n6396), .C(n7259), .Z(n7258) );
  HS65_LLS_XNOR2X6 U18609 ( .A(w1[0]), .B(n3006), .Z(n7259) );
  HS65_LL_OAI22X6 U18610 ( .A(n4071), .B(n9134), .C(n9126), .D(n4072), .Z(N34)
         );
  HS65_LLS_XNOR2X6 U18611 ( .A(w3[0]), .B(text_in_r[0]), .Z(n4071) );
  HS65_LLS_XOR3X2 U18612 ( .A(n2677), .B(n3218), .C(n4073), .Z(n4072) );
  HS65_LLS_XNOR2X6 U18613 ( .A(w3[0]), .B(n2674), .Z(n4073) );
  HS65_LL_OAI22X6 U18614 ( .A(n7563), .B(n9132), .C(n9128), .D(n7564), .Z(N137) );
  HS65_LLS_XNOR2X6 U18615 ( .A(w2[23]), .B(text_in_r[55]), .Z(n7563) );
  HS65_LLS_XOR3X2 U18616 ( .A(n7532), .B(n7535), .C(n7565), .Z(n7564) );
  HS65_LLS_XNOR2X6 U18617 ( .A(w2[23]), .B(n316), .Z(n7565) );
  HS65_LL_OAI22X6 U18618 ( .A(n2675), .B(n9131), .C(n9128), .D(n2676), .Z(N82)
         );
  HS65_LLS_XNOR2X6 U18619 ( .A(w3[24]), .B(text_in_r[24]), .Z(n2675) );
  HS65_LLS_XOR3X2 U18620 ( .A(n2654), .B(n2677), .C(n2678), .Z(n2676) );
  HS65_LLS_XNOR2X6 U18621 ( .A(w3[24]), .B(n183), .Z(n2678) );
  HS65_LL_OAI22X6 U18622 ( .A(n7541), .B(n9135), .C(n9122), .D(n7542), .Z(N150) );
  HS65_LLS_XNOR2X6 U18623 ( .A(w2[28]), .B(text_in_r[60]), .Z(n7541) );
  HS65_LLS_XOR3X2 U18624 ( .A(n7543), .B(n7544), .C(n7545), .Z(n7542) );
  HS65_LLS_XOR3X2 U18625 ( .A(n930), .B(n2754), .C(n2801), .Z(n7545) );
  HS65_LL_OAI22X6 U18626 ( .A(n5989), .B(n9130), .C(n9124), .D(n5990), .Z(N197) );
  HS65_LLS_XNOR2X6 U18627 ( .A(w1[19]), .B(text_in_r[83]), .Z(n5989) );
  HS65_LLS_XOR3X2 U18628 ( .A(n5986), .B(n5991), .C(n5992), .Z(n5990) );
  HS65_LLS_XOR3X2 U18629 ( .A(w1[19]), .B(n5962), .C(n2785), .Z(n5991) );
  HS65_LL_OAI22X6 U18630 ( .A(n7574), .B(n9132), .C(n9126), .D(n7575), .Z(N134) );
  HS65_LLS_XNOR2X6 U18631 ( .A(w2[20]), .B(text_in_r[52]), .Z(n7574) );
  HS65_LLS_XOR3X2 U18632 ( .A(n7576), .B(n7577), .C(n7578), .Z(n7575) );
  HS65_LLS_XOR3X2 U18633 ( .A(w2[20]), .B(n94), .C(n2778), .Z(n7577) );
  HS65_LL_OAI22X6 U18634 ( .A(n2693), .B(n9131), .C(n9128), .D(n2694), .Z(N70)
         );
  HS65_LLS_XNOR2X6 U18635 ( .A(w3[20]), .B(text_in_r[20]), .Z(n2693) );
  HS65_LLS_XOR3X2 U18636 ( .A(n2695), .B(n2696), .C(n2697), .Z(n2694) );
  HS65_LLS_XOR3X2 U18637 ( .A(n876), .B(n2660), .C(n2698), .Z(n2696) );
  HS65_LL_OAI22X6 U18638 ( .A(n4514), .B(n9135), .C(n9125), .D(n4515), .Z(N232) );
  HS65_LLS_XNOR2X6 U18639 ( .A(w0[6]), .B(text_in_r[102]), .Z(n4514) );
  HS65_LLS_XOR3X2 U18640 ( .A(n4351), .B(n4389), .C(n4516), .Z(n4515) );
  HS65_LLS_XNOR2X6 U18641 ( .A(w0[6]), .B(n3532), .Z(n4516) );
  HS65_LL_OAI22X6 U18642 ( .A(n6107), .B(n9129), .C(n9123), .D(n6108), .Z(N168) );
  HS65_LLS_XNOR2X6 U18643 ( .A(w1[6]), .B(text_in_r[70]), .Z(n6107) );
  HS65_LLS_XOR3X2 U18644 ( .A(n5944), .B(n5982), .C(n6109), .Z(n6108) );
  HS65_LLS_XNOR2X6 U18645 ( .A(w1[6]), .B(n3207), .Z(n6109) );
  HS65_LL_OAI22X6 U18646 ( .A(n2614), .B(n9132), .C(n9123), .D(n2615), .Z(N99)
         );
  HS65_LLS_XNOR2X6 U18647 ( .A(w2[1]), .B(text_in_r[33]), .Z(n2614) );
  HS65_LLS_XOR3X2 U18648 ( .A(n2616), .B(n2617), .C(n2618), .Z(n2615) );
  HS65_LLS_XOR3X2 U18649 ( .A(w2[1]), .B(n2619), .C(n2620), .Z(n2617) );
  HS65_LL_OAI22X6 U18650 ( .A(n5997), .B(n9129), .C(n9123), .D(n5998), .Z(N195) );
  HS65_LLS_XNOR2X6 U18651 ( .A(w1[17]), .B(text_in_r[81]), .Z(n5997) );
  HS65_LLS_XOR3X2 U18652 ( .A(n5986), .B(n5999), .C(n6000), .Z(n5998) );
  HS65_LLS_XOR3X2 U18653 ( .A(w1[17]), .B(n5971), .C(n2783), .Z(n5999) );
  HS65_LL_OAI22X6 U18654 ( .A(n4404), .B(n9134), .C(n9125), .D(n4405), .Z(N259) );
  HS65_LLS_XNOR2X6 U18655 ( .A(w0[17]), .B(text_in_r[113]), .Z(n4404) );
  HS65_LLS_XOR3X2 U18656 ( .A(n4393), .B(n4406), .C(n4407), .Z(n4405) );
  HS65_LLS_XOR3X2 U18657 ( .A(w0[17]), .B(n4378), .C(n2791), .Z(n4406) );
  HS65_LL_OAI22X6 U18658 ( .A(n2822), .B(n9136), .C(n9127), .D(n2823), .Z(N41)
         );
  HS65_LLS_XNOR2X6 U18659 ( .A(w3[7]), .B(text_in_r[7]), .Z(n2822) );
  HS65_LLS_XOR3X2 U18660 ( .A(n2654), .B(n2685), .C(n2824), .Z(n2823) );
  HS65_LLS_XNOR2X6 U18661 ( .A(w3[7]), .B(n404), .Z(n2824) );
  HS65_LL_OAI22X6 U18662 ( .A(n6018), .B(n9129), .C(n9123), .D(n6019), .Z(N181) );
  HS65_LLS_XNOR2X6 U18663 ( .A(w1[11]), .B(text_in_r[75]), .Z(n6018) );
  HS65_LLS_XOR3X2 U18664 ( .A(n6020), .B(n5992), .C(n6021), .Z(n6019) );
  HS65_LLS_XOR3X2 U18665 ( .A(w1[11]), .B(n2760), .C(n2784), .Z(n6021) );
  HS65_LL_OAI22X6 U18666 ( .A(n7603), .B(n9136), .C(n9127), .D(n7604), .Z(N118) );
  HS65_LLS_XNOR2X6 U18667 ( .A(w2[12]), .B(text_in_r[44]), .Z(n7603) );
  HS65_LLS_XOR3X2 U18668 ( .A(n7605), .B(n7578), .C(n7606), .Z(n7604) );
  HS65_LLS_XOR3X2 U18669 ( .A(w2[12]), .B(n2753), .C(n573), .Z(n7606) );
  HS65_LL_OAI22X6 U18670 ( .A(n7579), .B(n9132), .C(n9125), .D(n7580), .Z(N133) );
  HS65_LLS_XNOR2X6 U18671 ( .A(w2[19]), .B(text_in_r[51]), .Z(n7579) );
  HS65_LLS_XOR3X2 U18672 ( .A(n7576), .B(n7581), .C(n7582), .Z(n7580) );
  HS65_LLS_XOR3X2 U18673 ( .A(w2[19]), .B(n7555), .C(n2777), .Z(n7581) );
  HS65_LL_OAI22X6 U18674 ( .A(n4425), .B(n9135), .C(n9124), .D(n4426), .Z(N245) );
  HS65_LLS_XNOR2X6 U18675 ( .A(w0[11]), .B(text_in_r[107]), .Z(n4425) );
  HS65_LLS_XOR3X2 U18676 ( .A(n4427), .B(n4399), .C(n4428), .Z(n4426) );
  HS65_LLS_XOR3X2 U18677 ( .A(w0[11]), .B(n2768), .C(n2792), .Z(n4428) );
  HS65_LL_OAI22X6 U18678 ( .A(n5480), .B(n9130), .C(n9125), .D(n5481), .Z(N228) );
  HS65_LLS_XNOR2X6 U18679 ( .A(w0[2]), .B(text_in_r[98]), .Z(n5480) );
  HS65_LLS_XOR3X2 U18680 ( .A(n4369), .B(n4407), .C(n5482), .Z(n5481) );
  HS65_LLS_XNOR2X6 U18681 ( .A(w0[2]), .B(n3211), .Z(n5482) );
  HS65_LL_OAI22X6 U18682 ( .A(n7547), .B(n9136), .C(n9122), .D(n7548), .Z(N149) );
  HS65_LLS_XNOR2X6 U18683 ( .A(w2[27]), .B(text_in_r[59]), .Z(n7547) );
  HS65_LLS_XOR3X2 U18684 ( .A(n7549), .B(n7550), .C(n7551), .Z(n7548) );
  HS65_LLS_XOR3X2 U18685 ( .A(w2[27]), .B(n2753), .C(n2800), .Z(n7551) );
  HS65_LL_OAI22X6 U18686 ( .A(n7607), .B(n9132), .C(n9124), .D(n7608), .Z(N117) );
  HS65_LLS_XNOR2X6 U18687 ( .A(w2[11]), .B(text_in_r[43]), .Z(n7607) );
  HS65_LLS_XOR3X2 U18688 ( .A(n7609), .B(n7582), .C(n7610), .Z(n7608) );
  HS65_LLS_XOR3X2 U18689 ( .A(w2[11]), .B(n2752), .C(n2776), .Z(n7610) );
  HS65_LL_OAI22X6 U18690 ( .A(n4344), .B(n9135), .C(n9126), .D(n4345), .Z(N281) );
  HS65_LLS_XNOR2X6 U18691 ( .A(w0[31]), .B(text_in_r[127]), .Z(n4344) );
  HS65_LLS_XOR3X2 U18692 ( .A(n3532), .B(n4346), .C(n4347), .Z(n4345) );
  HS65_LLS_XOR3X2 U18693 ( .A(n2820), .B(n962), .C(n448), .Z(n4346) );
  HS65_LL_OAI22X6 U18694 ( .A(n5937), .B(n9130), .C(n9125), .D(n5938), .Z(N217) );
  HS65_LLS_XNOR2X6 U18695 ( .A(w1[31]), .B(text_in_r[95]), .Z(n5937) );
  HS65_LLS_XOR3X2 U18696 ( .A(n3207), .B(n5939), .C(n5940), .Z(n5938) );
  HS65_LLS_XOR3X2 U18697 ( .A(n2812), .B(n942), .C(n273), .Z(n5939) );
  HS65_LL_OAI22X6 U18698 ( .A(n5959), .B(n9130), .C(n9124), .D(n5960), .Z(N212) );
  HS65_LLS_XNOR2X6 U18699 ( .A(w1[26]), .B(text_in_r[90]), .Z(n5959) );
  HS65_LLS_XNOR3X2 U18700 ( .A(n3007), .B(n5961), .C(n5962), .Z(n5960) );
  HS65_LLS_XOR3X2 U18701 ( .A(n2760), .B(n939), .C(n2807), .Z(n5961) );
  HS65_LL_OAI22X6 U18702 ( .A(n5941), .B(n9130), .C(n9125), .D(n5942), .Z(N216) );
  HS65_LLS_XNOR2X6 U18703 ( .A(w1[30]), .B(text_in_r[94]), .Z(n5941) );
  HS65_LLS_XNOR3X2 U18704 ( .A(n3206), .B(n5943), .C(n5944), .Z(n5942) );
  HS65_LLS_XOR3X2 U18705 ( .A(n2764), .B(n941), .C(n2811), .Z(n5943) );
  HS65_LL_OAI22X6 U18706 ( .A(n4348), .B(n9136), .C(n9126), .D(n4349), .Z(N280) );
  HS65_LLS_XNOR2X6 U18707 ( .A(w0[30]), .B(text_in_r[126]), .Z(n4348) );
  HS65_LLS_XNOR3X2 U18708 ( .A(n3214), .B(n4350), .C(n4351), .Z(n4349) );
  HS65_LLS_XOR3X2 U18709 ( .A(n2772), .B(n961), .C(n2819), .Z(n4350) );
  HS65_LL_OAI22X6 U18710 ( .A(n4366), .B(n9136), .C(n9126), .D(n4367), .Z(N276) );
  HS65_LLS_XNOR2X6 U18711 ( .A(w0[26]), .B(text_in_r[122]), .Z(n4366) );
  HS65_LLS_XNOR3X2 U18712 ( .A(n3210), .B(n4368), .C(n4369), .Z(n4367) );
  HS65_LLS_XOR3X2 U18713 ( .A(n2768), .B(n958), .C(n2815), .Z(n4368) );
  HS65_LL_OAI22X6 U18714 ( .A(n4432), .B(n9133), .C(n9125), .D(n4433), .Z(N243) );
  HS65_LLS_XNOR2X6 U18715 ( .A(w0[9]), .B(text_in_r[105]), .Z(n4432) );
  HS65_LLS_XOR3X2 U18716 ( .A(n4407), .B(n4434), .C(n4435), .Z(n4433) );
  HS65_LLS_XOR3X2 U18717 ( .A(n2766), .B(w0[9]), .C(n2790), .Z(n4435) );
  HS65_LL_OAI22X6 U18718 ( .A(n7611), .B(n9132), .C(n9123), .D(n7612), .Z(N116) );
  HS65_LLS_XNOR2X6 U18719 ( .A(w2[10]), .B(text_in_r[42]), .Z(n7611) );
  HS65_LLS_XOR3X2 U18720 ( .A(n2800), .B(n7613), .C(n314), .Z(n7612) );
  HS65_LL_IVX9 U18721 ( .A(n7585), .Z(n314) );
  HS65_LL_OAI22X6 U18722 ( .A(n6022), .B(n9129), .C(n9123), .D(n6023), .Z(N180) );
  HS65_LLS_XNOR2X6 U18723 ( .A(w1[10]), .B(text_in_r[74]), .Z(n6022) );
  HS65_LLS_XNOR3X2 U18724 ( .A(n2808), .B(n6024), .C(n5995), .Z(n6023) );
  HS65_LLS_XOR3X2 U18725 ( .A(n2759), .B(n933), .C(n51), .Z(n6024) );
  HS65_LL_OAI22X6 U18726 ( .A(n7533), .B(n9130), .C(n9122), .D(n7534), .Z(N152) );
  HS65_LLS_XNOR2X6 U18727 ( .A(w2[30]), .B(text_in_r[62]), .Z(n7533) );
  HS65_LLS_XOR3X2 U18728 ( .A(n3003), .B(n7535), .C(n7536), .Z(n7534) );
  HS65_LLS_XOR3X2 U18729 ( .A(n2756), .B(n931), .C(n2803), .Z(n7536) );
  HS65_LL_AO22X9 U18730 ( .A(key[125]), .B(n9141), .C(n979), .D(n9118), .Z(
        \u0/N71 ) );
  HS65_LL_AO22X9 U18731 ( .A(key[103]), .B(n9140), .C(n1001), .D(n9118), .Z(
        \u0/N49 ) );
  HS65_LL_AO22X9 U18732 ( .A(key[15]), .B(n9121), .C(n1041), .D(n9146), .Z(
        \u0/N255 ) );
  HS65_LLS_XNOR2X6 U18733 ( .A(w3[15]), .B(n1042), .Z(n1041) );
  HS65_LL_AO22X9 U18734 ( .A(key[25]), .B(n9140), .C(n1021), .D(n9149), .Z(
        \u0/N265 ) );
  HS65_LLS_XNOR2X6 U18735 ( .A(w3[25]), .B(n1022), .Z(n1021) );
  HS65_LL_AO22X9 U18736 ( .A(key[22]), .B(ld), .C(n1027), .D(n9118), .Z(
        \u0/N262 ) );
  HS65_LLS_XNOR2X6 U18737 ( .A(w3[22]), .B(n1028), .Z(n1027) );
  HS65_LL_AO22X9 U18738 ( .A(key[6]), .B(ld), .C(n1059), .D(n9146), .Z(
        \u0/N246 ) );
  HS65_LLS_XNOR2X6 U18739 ( .A(w3[6]), .B(n1060), .Z(n1059) );
  HS65_LL_AO22X9 U18740 ( .A(key[2]), .B(ld), .C(n1067), .D(n9146), .Z(
        \u0/N242 ) );
  HS65_LLS_XNOR2X6 U18741 ( .A(w3[2]), .B(n1068), .Z(n1067) );
  HS65_LL_AO22X9 U18742 ( .A(key[18]), .B(ld), .C(n1035), .D(n9146), .Z(
        \u0/N258 ) );
  HS65_LLS_XNOR2X6 U18743 ( .A(w3[18]), .B(n1036), .Z(n1035) );
  HS65_LL_AO22X9 U18744 ( .A(key[0]), .B(n9140), .C(n1071), .D(n9147), .Z(
        \u0/N240 ) );
  HS65_LLS_XNOR2X6 U18745 ( .A(w3[0]), .B(n1072), .Z(n1071) );
  HS65_LL_AO22X9 U18746 ( .A(key[5]), .B(ld), .C(n1061), .D(n9146), .Z(
        \u0/N245 ) );
  HS65_LLS_XNOR2X6 U18747 ( .A(w3[5]), .B(n1062), .Z(n1061) );
  HS65_LL_AO22X9 U18748 ( .A(key[21]), .B(ld), .C(n1029), .D(n9148), .Z(
        \u0/N261 ) );
  HS65_LLS_XNOR2X6 U18749 ( .A(w3[21]), .B(n1030), .Z(n1029) );
  HS65_LL_AO22X9 U18750 ( .A(key[98]), .B(n9141), .C(n1006), .D(n9118), .Z(
        \u0/N44 ) );
  HS65_LL_AO22X9 U18751 ( .A(key[119]), .B(n9141), .C(n985), .D(n9144), .Z(
        \u0/N65 ) );
  HS65_LL_AO22X9 U18752 ( .A(key[67]), .B(n9142), .C(n1101), .D(n9144), .Z(
        \u0/N111 ) );
  HS65_LL_AO22X9 U18753 ( .A(key[91]), .B(n9141), .C(n1077), .D(n9147), .Z(
        \u0/N135 ) );
  HS65_LL_AO22X9 U18754 ( .A(key[81]), .B(n9142), .C(n1087), .D(n9147), .Z(
        \u0/N125 ) );
  HS65_LL_AO22X9 U18755 ( .A(key[83]), .B(n9141), .C(n1085), .D(n9147), .Z(
        \u0/N127 ) );
  HS65_LL_AO22X9 U18756 ( .A(key[80]), .B(n9142), .C(n1088), .D(n9147), .Z(
        \u0/N124 ) );
  HS65_LL_AO22X9 U18757 ( .A(key[88]), .B(n9141), .C(n1080), .D(n9147), .Z(
        \u0/N132 ) );
  HS65_LL_AO22X9 U18758 ( .A(key[73]), .B(n9142), .C(n1095), .D(n9148), .Z(
        \u0/N117 ) );
  HS65_LL_AO22X9 U18759 ( .A(key[78]), .B(n9142), .C(n1090), .D(n9147), .Z(
        \u0/N122 ) );
  HS65_LL_AO22X9 U18760 ( .A(key[65]), .B(n9142), .C(n1103), .D(n9144), .Z(
        \u0/N109 ) );
  HS65_LL_AO22X9 U18761 ( .A(key[75]), .B(n9142), .C(n1093), .D(n9144), .Z(
        \u0/N119 ) );
  HS65_LL_AO22X9 U18762 ( .A(key[64]), .B(n9142), .C(n1104), .D(n9149), .Z(
        \u0/N108 ) );
  HS65_LL_AO22X9 U18763 ( .A(key[72]), .B(n9142), .C(n1096), .D(n9144), .Z(
        \u0/N116 ) );
  HS65_LL_AO22X9 U18764 ( .A(key[70]), .B(n9142), .C(n1098), .D(n9148), .Z(
        \u0/N114 ) );
  HS65_LL_AO22X9 U18765 ( .A(key[86]), .B(n9141), .C(n1082), .D(n9147), .Z(
        \u0/N130 ) );
  HS65_LL_AO22X9 U18766 ( .A(key[31]), .B(n9140), .C(n1009), .D(n9149), .Z(
        \u0/N271 ) );
  HS65_LLS_XNOR2X6 U18767 ( .A(w3[31]), .B(n1010), .Z(n1009) );
  HS65_LL_AO22X9 U18768 ( .A(key[12]), .B(ld), .C(n1047), .D(n9146), .Z(
        \u0/N252 ) );
  HS65_LLS_XNOR2X6 U18769 ( .A(w3[12]), .B(n1048), .Z(n1047) );
  HS65_LL_AO22X9 U18770 ( .A(key[24]), .B(n9140), .C(n1023), .D(n9149), .Z(
        \u0/N264 ) );
  HS65_LLS_XNOR2X6 U18771 ( .A(w3[24]), .B(n1024), .Z(n1023) );
  HS65_LL_AO22X9 U18772 ( .A(key[16]), .B(ld), .C(n1039), .D(n9146), .Z(
        \u0/N256 ) );
  HS65_LLS_XNOR2X6 U18773 ( .A(w3[16]), .B(n1040), .Z(n1039) );
  HS65_LL_AO22X9 U18774 ( .A(key[8]), .B(n9141), .C(n1055), .D(n9146), .Z(
        \u0/N248 ) );
  HS65_LLS_XNOR2X6 U18775 ( .A(w3[8]), .B(n1056), .Z(n1055) );
  HS65_LL_AO22X9 U18776 ( .A(key[20]), .B(n9140), .C(n1031), .D(n9149), .Z(
        \u0/N260 ) );
  HS65_LLS_XNOR2X6 U18777 ( .A(w3[20]), .B(n1032), .Z(n1031) );
  HS65_LL_AO22X9 U18778 ( .A(key[1]), .B(ld), .C(n1069), .D(n9146), .Z(
        \u0/N241 ) );
  HS65_LLS_XNOR2X6 U18779 ( .A(w3[1]), .B(n1070), .Z(n1069) );
  HS65_LL_AO22X9 U18780 ( .A(key[7]), .B(ld), .C(n1057), .D(n9146), .Z(
        \u0/N247 ) );
  HS65_LLS_XNOR2X6 U18781 ( .A(w3[7]), .B(n1058), .Z(n1057) );
  HS65_LL_AO22X9 U18782 ( .A(key[23]), .B(n9140), .C(n1025), .D(n9149), .Z(
        \u0/N263 ) );
  HS65_LLS_XNOR2X6 U18783 ( .A(w3[23]), .B(n1026), .Z(n1025) );
  HS65_LL_AO22X9 U18784 ( .A(key[19]), .B(ld), .C(n1033), .D(n9146), .Z(
        \u0/N259 ) );
  HS65_LLS_XNOR2X6 U18785 ( .A(w3[19]), .B(n1034), .Z(n1033) );
  HS65_LL_AO22X9 U18786 ( .A(key[17]), .B(ld), .C(n1037), .D(n9146), .Z(
        \u0/N257 ) );
  HS65_LLS_XNOR2X6 U18787 ( .A(w3[17]), .B(n1038), .Z(n1037) );
  HS65_LL_AO22X9 U18788 ( .A(key[3]), .B(ld), .C(n1065), .D(n9146), .Z(
        \u0/N243 ) );
  HS65_LLS_XNOR2X6 U18789 ( .A(w3[3]), .B(n1066), .Z(n1065) );
  HS65_LL_AO22X9 U18790 ( .A(key[77]), .B(n9142), .C(n1091), .D(n9147), .Z(
        \u0/N121 ) );
  HS65_LL_AO22X9 U18791 ( .A(key[93]), .B(n9141), .C(n1075), .D(n9147), .Z(
        \u0/N137 ) );
  HS65_LL_AO22X9 U18792 ( .A(key[71]), .B(n9142), .C(n1097), .D(n9144), .Z(
        \u0/N115 ) );
  HS65_LL_AO22X9 U18793 ( .A(key[14]), .B(ld), .C(n1043), .D(n9146), .Z(
        \u0/N254 ) );
  HS65_LLS_XNOR2X6 U18794 ( .A(w3[14]), .B(n1044), .Z(n1043) );
  HS65_LL_AO22X9 U18795 ( .A(key[30]), .B(n9140), .C(n1011), .D(n9149), .Z(
        \u0/N270 ) );
  HS65_LLS_XNOR2X6 U18796 ( .A(w3[30]), .B(n1012), .Z(n1011) );
  HS65_LL_AO22X9 U18797 ( .A(key[10]), .B(ld), .C(n1051), .D(n9146), .Z(
        \u0/N250 ) );
  HS65_LLS_XNOR2X6 U18798 ( .A(w3[10]), .B(n1052), .Z(n1051) );
  HS65_LL_AO22X9 U18799 ( .A(key[13]), .B(ld), .C(n1045), .D(n9146), .Z(
        \u0/N253 ) );
  HS65_LLS_XNOR2X6 U18800 ( .A(w3[13]), .B(n1046), .Z(n1045) );
  HS65_LL_AO22X9 U18801 ( .A(key[68]), .B(n9142), .C(n1100), .D(n9144), .Z(
        \u0/N112 ) );
  HS65_LL_AO22X9 U18802 ( .A(key[76]), .B(n9142), .C(n1092), .D(n9148), .Z(
        \u0/N120 ) );
  HS65_LL_AO22X9 U18803 ( .A(key[87]), .B(n9141), .C(n1081), .D(n9147), .Z(
        \u0/N131 ) );
  HS65_LL_AO22X9 U18804 ( .A(key[66]), .B(n9142), .C(n1102), .D(n9144), .Z(
        \u0/N110 ) );
  HS65_LL_AO22X9 U18805 ( .A(key[92]), .B(n9141), .C(n1076), .D(n9147), .Z(
        \u0/N136 ) );
  HS65_LL_AO22X9 U18806 ( .A(key[84]), .B(n9141), .C(n1084), .D(n9147), .Z(
        \u0/N128 ) );
  HS65_LL_AO22X9 U18807 ( .A(key[82]), .B(n9141), .C(n1086), .D(n9147), .Z(
        \u0/N126 ) );
  HS65_LL_AO22X9 U18808 ( .A(key[85]), .B(n9141), .C(n1083), .D(n9147), .Z(
        \u0/N129 ) );
  HS65_LL_AO22X9 U18809 ( .A(key[69]), .B(n9142), .C(n1099), .D(n9148), .Z(
        \u0/N113 ) );
  HS65_LL_AO22X9 U18810 ( .A(key[95]), .B(n9141), .C(n1073), .D(n9147), .Z(
        \u0/N139 ) );
  HS65_LL_AO22X9 U18811 ( .A(key[74]), .B(n9142), .C(n1094), .D(n9144), .Z(
        \u0/N118 ) );
  HS65_LL_AO22X9 U18812 ( .A(key[79]), .B(n9142), .C(n1089), .D(n9147), .Z(
        \u0/N123 ) );
  HS65_LL_AO22X9 U18813 ( .A(key[90]), .B(n9141), .C(n1078), .D(n9147), .Z(
        \u0/N134 ) );
  HS65_LL_AO22X9 U18814 ( .A(key[111]), .B(n9140), .C(n993), .D(n9144), .Z(
        \u0/N57 ) );
  HS65_LL_AO22X9 U18815 ( .A(key[106]), .B(n9140), .C(n998), .D(n9149), .Z(
        \u0/N52 ) );
  HS65_LL_AO22X9 U18816 ( .A(key[122]), .B(n9142), .C(n982), .D(n9144), .Z(
        \u0/N68 ) );
  HS65_LL_AO22X9 U18817 ( .A(n9116), .B(key[127]), .C(n977), .D(n9148), .Z(
        \u0/N73 ) );
  HS65_LL_AO22X9 U18818 ( .A(key[114]), .B(n9140), .C(n990), .D(n9149), .Z(
        \u0/N60 ) );
  HS65_LL_AO22X9 U18819 ( .A(key[89]), .B(n9141), .C(n1079), .D(n9147), .Z(
        \u0/N133 ) );
  HS65_LL_AO22X9 U18820 ( .A(key[94]), .B(n9141), .C(n1074), .D(n9147), .Z(
        \u0/N138 ) );
  HS65_LL_IVX9 U18821 ( .A(\u0/r0/rcnt [0]), .Z(n964) );
  HS65_LL_NOR2X6 U18822 ( .A(sa00[3]), .B(sa00[2]), .Z(n5809) );
  HS65_LL_OAI22X6 U18823 ( .A(n2726), .B(n9131), .C(n9127), .D(n2727), .Z(N55)
         );
  HS65_LLS_XNOR2X6 U18824 ( .A(w3[13]), .B(text_in_r[13]), .Z(n2726) );
  HS65_LLS_XNOR3X2 U18825 ( .A(n2698), .B(n2728), .C(n2690), .Z(n2727) );
  HS65_LLS_XOR3X2 U18826 ( .A(n2634), .B(n836), .C(n187), .Z(n2728) );
  HS65_LL_OAI22X6 U18827 ( .A(n5945), .B(n9130), .C(n9124), .D(n5946), .Z(N215) );
  HS65_LLS_XNOR2X6 U18828 ( .A(w1[29]), .B(text_in_r[93]), .Z(n5945) );
  HS65_LLS_XNOR3X2 U18829 ( .A(n3205), .B(n5947), .C(n5948), .Z(n5946) );
  HS65_LLS_XOR3X2 U18830 ( .A(n2763), .B(w1[29]), .C(n2810), .Z(n5947) );
  HS65_LL_OAI22X6 U18831 ( .A(n4352), .B(n9136), .C(n9126), .D(n4353), .Z(N279) );
  HS65_LLS_XNOR2X6 U18832 ( .A(w0[29]), .B(text_in_r[125]), .Z(n4352) );
  HS65_LLS_XNOR3X2 U18833 ( .A(n3213), .B(n4354), .C(n4355), .Z(n4353) );
  HS65_LLS_XOR3X2 U18834 ( .A(n2771), .B(w0[29]), .C(n2818), .Z(n4354) );
  HS65_LL_NOR3X4 U18835 ( .A(dcnt[1]), .B(dcnt[2]), .C(dcnt[0]), .Z(n2612) );
  HS65_LLS_XOR2X6 U18836 ( .A(\u0/r0/rcnt [1]), .B(n964), .Z(n968) );
  HS65_LLS_XOR2X6 U18837 ( .A(n975), .B(\u0/r0/rcnt [3]), .Z(n966) );
  HS65_LL_NAND2X7 U18838 ( .A(\u0/r0/rcnt [2]), .B(n976), .Z(n975) );
  HS65_LL_NAND2X7 U18839 ( .A(n974), .B(\u0/r0/rcnt [0]), .Z(n973) );
  HS65_LL_OAI32X5 U18840 ( .A(n706), .B(\u0/r0/rcnt [0]), .C(n972), .D(n9139), 
        .E(n973), .Z(\u0/r0/N73 ) );
  HS65_LLS_XNOR2X6 U18841 ( .A(n976), .B(\u0/r0/rcnt [2]), .Z(n971) );
  HS65_LLS_XNOR2X6 U18842 ( .A(n2749), .B(w3[15]), .Z(N466) );
  HS65_LLS_XNOR2X6 U18843 ( .A(n2896), .B(w3[25]), .Z(N408) );
  HS65_LLS_XNOR2X6 U18844 ( .A(n2659), .B(w3[18]), .Z(N439) );
  HS65_LLS_XNOR2X6 U18845 ( .A(n2637), .B(w3[6]), .Z(N499) );
  HS65_LLS_XNOR2X6 U18846 ( .A(n2745), .B(w3[0]), .Z(N505) );
  HS65_LLS_XNOR2X6 U18847 ( .A(n2627), .B(w3[22]), .Z(N435) );
  HS65_LLS_XNOR2X6 U18848 ( .A(n2666), .B(w3[2]), .Z(N503) );
  HS65_LLS_XNOR2X6 U18849 ( .A(n2634), .B(w3[21]), .Z(N436) );
  HS65_LLS_XNOR2X6 U18850 ( .A(n2644), .B(w3[5]), .Z(N500) );
  HS65_LL_AOI112X4 U18851 ( .A(n2), .B(n2612), .C(N0), .D(n9137), .Z(n2610) );
  HS65_LLS_XNOR2X6 U18852 ( .A(n2651), .B(w3[4]), .Z(N501) );
  HS65_LLS_XNOR2X6 U18853 ( .A(n2897), .B(w3[26]), .Z(N407) );
  HS65_LLS_XNOR2X6 U18854 ( .A(n2641), .B(w3[20]), .Z(N437) );
  HS65_LLS_XNOR2X6 U18855 ( .A(n2663), .B(w3[17]), .Z(N440) );
  HS65_LLS_XNOR2X6 U18856 ( .A(n2653), .B(w3[19]), .Z(N438) );
  HS65_LLS_XNOR2X6 U18857 ( .A(n2733), .B(w3[3]), .Z(N502) );
  HS65_LL_AND2X4 U18858 ( .A(sa00[7]), .B(sa00[6]), .Z(n5801) );
  HS65_LL_IVX9 U18859 ( .A(w1[25]), .Z(n938) );
  HS65_LL_IVX9 U18860 ( .A(w1[30]), .Z(n941) );
  HS65_LL_IVX9 U18861 ( .A(w0[3]), .Z(n944) );
  HS65_LL_OAI31X5 U18862 ( .A(n963), .B(\u0/r0/rcnt [0]), .C(n967), .D(n969), 
        .Z(\u0/r0/N75 ) );
  HS65_LL_IVX9 U18863 ( .A(w0[15]), .Z(n949) );
  HS65_LL_IVX9 U18864 ( .A(w0[10]), .Z(n947) );
  HS65_LL_NOR2X6 U18865 ( .A(n9139), .B(\u0/r0/rcnt [0]), .Z(\u0/r0/N78 ) );
  HS65_LLS_XNOR2X6 U18866 ( .A(n2898), .B(w2[24]), .Z(N401) );
  HS65_LLS_XNOR2X6 U18867 ( .A(n2804), .B(w2[22]), .Z(N427) );
  HS65_LLS_XNOR2X6 U18868 ( .A(n2755), .B(w2[5]), .Z(N492) );
  HS65_LLS_XNOR2X6 U18869 ( .A(n2762), .B(w1[4]), .Z(N485) );
  HS65_LL_IVX9 U18870 ( .A(w0[14]), .Z(n948) );
  HS65_LLS_XNOR2X6 U18871 ( .A(n2786), .B(w1[12]), .Z(N453) );
  HS65_LLS_XNOR2X6 U18872 ( .A(n2813), .B(w1[23]), .Z(N418) );
  HS65_LLS_XNOR2X6 U18873 ( .A(n2760), .B(w1[2]), .Z(N487) );
  HS65_LLS_XOR2X6 U18874 ( .A(n3206), .B(w1[29]), .Z(N388) );
  HS65_LLS_XOR2X6 U18875 ( .A(n2787), .B(w1[13]), .Z(N452) );
  HS65_LL_IVX9 U18876 ( .A(w0[30]), .Z(n961) );
  HS65_LL_IVX9 U18877 ( .A(w0[25]), .Z(n957) );
  HS65_LL_IVX9 U18878 ( .A(w0[1]), .Z(n943) );
  HS65_LLS_XOR2X6 U18879 ( .A(n2765), .B(w1[7]), .Z(N482) );
  HS65_LL_IVX9 U18880 ( .A(w0[17]), .Z(n951) );
  HS65_LL_IVX9 U18881 ( .A(w0[19]), .Z(n953) );
  HS65_LL_IVX9 U18882 ( .A(w0[16]), .Z(n950) );
  HS65_LL_IVX9 U18883 ( .A(w0[27]), .Z(n959) );
  HS65_LL_NOR2AX3 U18884 ( .A(\u0/r0/rcnt [1]), .B(n964), .Z(n976) );
  HS65_LL_IVX9 U18885 ( .A(w0[31]), .Z(n962) );
  HS65_LL_IVX9 U18886 ( .A(w0[26]), .Z(n958) );
  HS65_LLS_XNOR2X6 U18887 ( .A(n2791), .B(w0[9]), .Z(N448) );
  HS65_LLS_XNOR2X6 U18888 ( .A(n2783), .B(w1[9]), .Z(N456) );
  HS65_LLS_XNOR2X6 U18889 ( .A(n2779), .B(w2[13]), .Z(N460) );
  HS65_LLS_XNOR2X6 U18890 ( .A(n2780), .B(w2[14]), .Z(N459) );
  HS65_LLS_XNOR2X6 U18891 ( .A(n2788), .B(w1[14]), .Z(N451) );
  HS65_LLS_XNOR2X6 U18892 ( .A(n3005), .B(w2[31]), .Z(N394) );
  HS65_LLS_XNOR2X6 U18893 ( .A(n3003), .B(w2[29]), .Z(N396) );
  HS65_LL_IVX9 U18894 ( .A(w0[4]), .Z(n945) );
  HS65_LLS_XNOR2X6 U18895 ( .A(n2795), .B(w0[13]), .Z(N444) );
  HS65_LL_NOR3X4 U18896 ( .A(n967), .B(\u0/r0/rcnt [0]), .C(n968), .Z(
        \u0/r0/N77 ) );
  HS65_LL_IVX9 U18897 ( .A(dcnt[0]), .Z(n5) );
  HS65_LLS_XNOR2X6 U18898 ( .A(n2759), .B(w1[1]), .Z(N488) );
  HS65_LLS_XNOR2X6 U18899 ( .A(n2753), .B(w2[3]), .Z(N494) );
  HS65_LLS_XNOR2X6 U18900 ( .A(n2777), .B(w2[11]), .Z(N462) );
  HS65_LLS_XNOR2X6 U18901 ( .A(n2785), .B(w1[11]), .Z(N454) );
  HS65_LLS_XNOR2X6 U18902 ( .A(n2793), .B(w0[11]), .Z(N446) );
  HS65_LLS_XNOR2X6 U18903 ( .A(n2620), .B(w2[25]), .Z(N400) );
  HS65_LLS_XNOR2X6 U18904 ( .A(n2775), .B(w2[9]), .Z(N464) );
  HS65_LLS_XNOR2X6 U18905 ( .A(n2794), .B(w0[12]), .Z(N445) );
  HS65_LL_IVX9 U18906 ( .A(w0[20]), .Z(n954) );
  HS65_LL_IVX9 U18907 ( .A(w0[18]), .Z(n952) );
  HS65_LL_IVX9 U18908 ( .A(w0[21]), .Z(n955) );
  HS65_LL_IVX9 U18909 ( .A(w0[5]), .Z(n946) );
  HS65_LLS_XNOR2X6 U18910 ( .A(n2820), .B(w0[22]), .Z(N411) );
  HS65_LLS_XNOR2X6 U18911 ( .A(n2805), .B(w2[23]), .Z(N426) );
  HS65_LLS_XNOR2X6 U18912 ( .A(n2812), .B(w1[22]), .Z(N419) );
  HS65_LLS_XNOR2X6 U18913 ( .A(n2772), .B(w0[6]), .Z(N475) );
  HS65_LLS_XNOR2X6 U18914 ( .A(n2764), .B(w1[6]), .Z(N483) );
  HS65_LLS_XNOR2X6 U18915 ( .A(n2756), .B(w2[6]), .Z(N491) );
  HS65_LLS_XNOR2X6 U18916 ( .A(n2758), .B(w1[0]), .Z(N489) );
  HS65_LLS_XNOR2X6 U18917 ( .A(n2750), .B(w2[0]), .Z(N497) );
  HS65_LLS_XNOR2X6 U18918 ( .A(n2752), .B(w2[2]), .Z(N495) );
  HS65_LLS_XNOR2X6 U18919 ( .A(n2782), .B(w1[8]), .Z(N457) );
  HS65_LLS_XOR2X6 U18920 ( .A(n2776), .B(w2[10]), .Z(N463) );
  HS65_LLS_XNOR2X6 U18921 ( .A(n2821), .B(w0[23]), .Z(N410) );
  HS65_LLS_XNOR2X6 U18922 ( .A(n2768), .B(w0[2]), .Z(N479) );
  HS65_LLS_XOR2X6 U18923 ( .A(n3009), .B(w1[27]), .Z(N390) );
  HS65_LLS_XOR2X6 U18924 ( .A(n2754), .B(w2[4]), .Z(N493) );
  HS65_LLS_XOR2X6 U18925 ( .A(n2761), .B(w1[3]), .Z(N486) );
  HS65_LLS_XOR2X6 U18926 ( .A(n2778), .B(w2[12]), .Z(N461) );
  HS65_LLS_XOR2X6 U18927 ( .A(n2809), .B(w1[19]), .Z(N422) );
  HS65_LLS_XOR2X6 U18928 ( .A(n2807), .B(w1[17]), .Z(N424) );
  HS65_LLS_XOR2X6 U18929 ( .A(n2751), .B(w2[1]), .Z(N496) );
  HS65_LLS_XOR2X6 U18930 ( .A(n3214), .B(w0[29]), .Z(N380) );
  HS65_LLS_XOR2X6 U18931 ( .A(n2781), .B(w2[15]), .Z(N458) );
  HS65_LLS_XOR2X6 U18932 ( .A(n3006), .B(w1[24]), .Z(N393) );
  HS65_LLS_XOR2X6 U18933 ( .A(n2774), .B(w2[8]), .Z(N465) );
  HS65_LLS_XOR2X6 U18934 ( .A(n2766), .B(w0[0]), .Z(N481) );
  HS65_LLS_XOR2X6 U18935 ( .A(n2790), .B(w0[8]), .Z(N449) );
  HS65_LLS_XOR2X6 U18936 ( .A(n2806), .B(w1[16]), .Z(N425) );
  HS65_LLS_XOR2X6 U18937 ( .A(n2773), .B(w0[7]), .Z(N474) );
  HS65_LL_IVX9 U18938 ( .A(w1[26]), .Z(n939) );
  HS65_LL_IVX9 U18939 ( .A(w1[15]), .Z(n934) );
  HS65_LL_IVX9 U18940 ( .A(w1[10]), .Z(n933) );
  HS65_LL_IVX9 U18941 ( .A(w1[31]), .Z(n942) );
  HS65_LL_IVX9 U18942 ( .A(w2[30]), .Z(n931) );
  HS65_LL_IVX9 U18943 ( .A(w2[26]), .Z(n928) );
  HS65_LL_OAI22X6 U18944 ( .A(n2688), .B(n9131), .C(n9128), .D(n2689), .Z(N71)
         );
  HS65_LLS_XNOR2X6 U18945 ( .A(w3[21]), .B(text_in_r[21]), .Z(n2688) );
  HS65_LLS_XOR3X2 U18946 ( .A(n2649), .B(n2690), .C(n2691), .Z(n2689) );
  HS65_LLS_XNOR2X6 U18947 ( .A(w3[21]), .B(n2692), .Z(n2691) );
  HS65_LL_OAI22X6 U18948 ( .A(n3010), .B(n9136), .C(n9127), .D(n3011), .Z(N39)
         );
  HS65_LLS_XNOR2X6 U18949 ( .A(w3[5]), .B(text_in_r[5]), .Z(n3010) );
  HS65_LLS_XOR3X2 U18950 ( .A(n2643), .B(n2697), .C(n3012), .Z(n3011) );
  HS65_LLS_XNOR2X6 U18951 ( .A(w3[5]), .B(n2638), .Z(n3012) );
  HS65_LL_IVX9 U18952 ( .A(w0[24]), .Z(n956) );
  HS65_LL_IVX9 U18953 ( .A(w2[28]), .Z(n930) );
  HS65_LL_IVX9 U18954 ( .A(w0[28]), .Z(n960) );
  HS65_LL_OAI22X6 U18955 ( .A(n6204), .B(n9129), .C(n9122), .D(n6205), .Z(N167) );
  HS65_LLS_XNOR2X6 U18956 ( .A(w1[5]), .B(text_in_r[69]), .Z(n6204) );
  HS65_LLS_XOR3X2 U18957 ( .A(n5948), .B(n5988), .C(n6206), .Z(n6205) );
  HS65_LLS_XNOR2X6 U18958 ( .A(w1[5]), .B(n3206), .Z(n6206) );
  HS65_LL_OAI22X6 U18959 ( .A(n7600), .B(n9136), .C(n9128), .D(n7601), .Z(N119) );
  HS65_LLS_XNOR2X6 U18960 ( .A(w2[13]), .B(text_in_r[45]), .Z(n7600) );
  HS65_LLS_XNOR3X2 U18961 ( .A(n2803), .B(n7602), .C(n7572), .Z(n7601) );
  HS65_LLS_XOR3X2 U18962 ( .A(n2754), .B(w2[13]), .C(n2778), .Z(n7602) );
  HS65_LL_NOR3X4 U18963 ( .A(n5114), .B(dcnt[1]), .C(n5), .Z(N23) );
  HS65_LL_NAND3AX6 U18964 ( .A(dcnt[2]), .B(n2), .C(n9144), .Z(n5114) );
  HS65_LL_OAI22X6 U18965 ( .A(n7570), .B(n9132), .C(n9124), .D(n7571), .Z(N135) );
  HS65_LLS_XNOR2X6 U18966 ( .A(w2[21]), .B(text_in_r[53]), .Z(n7570) );
  HS65_LLS_XOR3X2 U18967 ( .A(n7544), .B(n7572), .C(n7573), .Z(n7571) );
  HS65_LLS_XNOR2X6 U18968 ( .A(w2[21]), .B(n572), .Z(n7573) );
  HS65_LLS_XNOR2X6 U18969 ( .A(n2796), .B(w0[14]), .Z(N443) );
  HS65_LLS_XNOR2X6 U18970 ( .A(n2767), .B(w0[1]), .Z(N480) );
  HS65_LLS_XNOR2X6 U18971 ( .A(n2770), .B(w0[4]), .Z(N477) );
  HS65_LL_OAI22X6 U18972 ( .A(n4611), .B(n9134), .C(n9125), .D(n4612), .Z(N231) );
  HS65_LLS_XNOR2X6 U18973 ( .A(w0[5]), .B(text_in_r[101]), .Z(n4611) );
  HS65_LLS_XOR3X2 U18974 ( .A(n4355), .B(n4395), .C(n4613), .Z(n4612) );
  HS65_LLS_XNOR2X6 U18975 ( .A(w0[5]), .B(n3214), .Z(n4613) );
  HS65_LL_OAI31X5 U18976 ( .A(n2), .B(n2612), .C(n1), .D(n705), .Z(n9113) );
  HS65_LL_OAI22X6 U18977 ( .A(n717), .B(n9145), .C(n994), .D(n9138), .Z(
        \u0/N56 ) );
  HS65_LL_IVX9 U18978 ( .A(key[110]), .Z(n717) );
  HS65_LL_OAI22X6 U18979 ( .A(n713), .B(n9145), .C(n986), .D(n9137), .Z(
        \u0/N64 ) );
  HS65_LL_IVX9 U18980 ( .A(key[118]), .Z(n713) );
  HS65_LL_OAI22X6 U18981 ( .A(n709), .B(n9145), .C(n978), .D(n9137), .Z(
        \u0/N72 ) );
  HS65_LL_IVX9 U18982 ( .A(key[126]), .Z(n709) );
  HS65_LL_OAI22X6 U18983 ( .A(n714), .B(n9145), .C(n989), .D(n9138), .Z(
        \u0/N61 ) );
  HS65_LL_IVX9 U18984 ( .A(key[115]), .Z(n714) );
  HS65_LL_OAI22X6 U18985 ( .A(n718), .B(n9145), .C(n997), .D(n9138), .Z(
        \u0/N53 ) );
  HS65_LL_IVX9 U18986 ( .A(key[107]), .Z(n718) );
  HS65_LL_OAI22X6 U18987 ( .A(n721), .B(n9145), .C(n1002), .D(n9138), .Z(
        \u0/N48 ) );
  HS65_LL_IVX9 U18988 ( .A(key[102]), .Z(n721) );
  HS65_LL_OAI22X6 U18989 ( .A(n715), .B(n9145), .C(n991), .D(n9138), .Z(
        \u0/N59 ) );
  HS65_LL_IVX9 U18990 ( .A(key[113]), .Z(n715) );
  HS65_LL_OAI22X6 U18991 ( .A(n710), .B(n9145), .C(n981), .D(n9137), .Z(
        \u0/N69 ) );
  HS65_LL_IVX9 U18992 ( .A(key[123]), .Z(n710) );
  HS65_LL_OAI22X6 U18993 ( .A(n719), .B(n9145), .C(n999), .D(n9138), .Z(
        \u0/N51 ) );
  HS65_LL_IVX9 U18994 ( .A(key[105]), .Z(n719) );
  HS65_LL_OAI22X6 U18995 ( .A(n711), .B(n9145), .C(n983), .D(n9137), .Z(
        \u0/N67 ) );
  HS65_LL_IVX9 U18996 ( .A(key[121]), .Z(n711) );
  HS65_LL_OAI22X6 U18997 ( .A(n712), .B(n9145), .C(n984), .D(n9137), .Z(
        \u0/N66 ) );
  HS65_LL_IVX9 U18998 ( .A(key[120]), .Z(n712) );
  HS65_LL_OAI22X6 U18999 ( .A(n716), .B(n9145), .C(n992), .D(n9138), .Z(
        \u0/N58 ) );
  HS65_LL_IVX9 U19000 ( .A(key[112]), .Z(n716) );
  HS65_LL_OAI22X6 U19001 ( .A(n720), .B(n9145), .C(n1000), .D(n9139), .Z(
        \u0/N50 ) );
  HS65_LL_IVX9 U19002 ( .A(key[104]), .Z(n720) );
  HS65_LL_OAI22X6 U19003 ( .A(n723), .B(n9149), .C(n1007), .D(n9139), .Z(
        \u0/N43 ) );
  HS65_LL_IVX9 U19004 ( .A(key[97]), .Z(n723) );
  HS65_LL_OAI22X6 U19005 ( .A(n722), .B(n9149), .C(n1005), .D(n9139), .Z(
        \u0/N45 ) );
  HS65_LL_IVX9 U19006 ( .A(key[99]), .Z(n722) );
  HS65_LL_OAI22X6 U19007 ( .A(n724), .B(n9143), .C(n1008), .D(n9139), .Z(
        \u0/N42 ) );
  HS65_LL_IVX9 U19008 ( .A(key[96]), .Z(n724) );
  HS65_LL_OAI21X3 U19009 ( .A(dcnt[0]), .B(n1), .C(n705), .Z(n9114) );
  HS65_LL_NOR2X6 U19010 ( .A(n9144), .B(N0), .Z(n2613) );
  HS65_LLS_XOR2X6 U19011 ( .A(n2757), .B(w2[7]), .Z(N490) );
  HS65_LLS_XOR2X6 U19012 ( .A(n3001), .B(w2[27]), .Z(N398) );
  HS65_LLS_XOR2X6 U19013 ( .A(n2802), .B(w2[20]), .Z(N429) );
  HS65_LLS_XOR2X6 U19014 ( .A(n2801), .B(w2[19]), .Z(N430) );
  HS65_LLS_XOR2X6 U19015 ( .A(n2763), .B(w1[5]), .Z(N484) );
  HS65_LLS_XOR2X6 U19016 ( .A(n2803), .B(w2[21]), .Z(N428) );
  HS65_LLS_XOR2X6 U19017 ( .A(n2811), .B(w1[21]), .Z(N420) );
  HS65_LLS_XOR2X6 U19018 ( .A(n2799), .B(w2[17]), .Z(N432) );
  HS65_LLS_XOR2X6 U19019 ( .A(n2808), .B(w1[18]), .Z(N423) );
  HS65_LLS_XOR2X6 U19020 ( .A(n2800), .B(w2[18]), .Z(N431) );
  HS65_LLS_XOR2X6 U19021 ( .A(n2798), .B(w2[16]), .Z(N433) );
  HS65_LL_OAI22X6 U19022 ( .A(n7537), .B(n9135), .C(n9122), .D(n7538), .Z(N151) );
  HS65_LLS_XNOR2X6 U19023 ( .A(w2[29]), .B(text_in_r[61]), .Z(n7537) );
  HS65_LLS_XNOR3X2 U19024 ( .A(n3002), .B(n7539), .C(n7540), .Z(n7538) );
  HS65_LLS_XOR3X2 U19025 ( .A(n361), .B(w2[29]), .C(n2802), .Z(n7539) );
  HS65_LLS_XOR2X6 U19026 ( .A(n3205), .B(w1[28]), .Z(N389) );
  HS65_LLS_XOR2X6 U19027 ( .A(n2810), .B(w1[20]), .Z(N421) );
  HS65_LL_OAI22X6 U19028 ( .A(n2639), .B(n9131), .C(n9128), .D(n2640), .Z(N87)
         );
  HS65_LLS_XNOR2X6 U19029 ( .A(w3[29]), .B(text_in_r[29]), .Z(n2639) );
  HS65_LLS_XOR3X2 U19030 ( .A(n2641), .B(n2642), .C(n2643), .Z(n2640) );
  HS65_LLS_XOR3X2 U19031 ( .A(n2644), .B(n918), .C(n2645), .Z(n2642) );
  HS65_LL_OAI22X6 U19032 ( .A(n5980), .B(n9130), .C(n9124), .D(n5981), .Z(N199) );
  HS65_LLS_XNOR2X6 U19033 ( .A(w1[21]), .B(text_in_r[85]), .Z(n5980) );
  HS65_LLS_XOR3X2 U19034 ( .A(n5952), .B(n5982), .C(n5983), .Z(n5981) );
  HS65_LLS_XNOR2X6 U19035 ( .A(w1[21]), .B(n2787), .Z(n5983) );
  HS65_LL_OAI22X6 U19036 ( .A(n4387), .B(n9135), .C(n9123), .D(n4388), .Z(N263) );
  HS65_LLS_XNOR2X6 U19037 ( .A(w0[21]), .B(text_in_r[117]), .Z(n4387) );
  HS65_LLS_XOR3X2 U19038 ( .A(n4359), .B(n4389), .C(n4390), .Z(n4388) );
  HS65_LLS_XNOR2X6 U19039 ( .A(w0[21]), .B(n230), .Z(n4390) );
  HS65_LL_OAI22X6 U19040 ( .A(n8020), .B(n9132), .C(n9122), .D(n8021), .Z(N103) );
  HS65_LLS_XNOR2X6 U19041 ( .A(w2[5]), .B(text_in_r[37]), .Z(n8020) );
  HS65_LLS_XOR3X2 U19042 ( .A(n7540), .B(n7578), .C(n8022), .Z(n8021) );
  HS65_LLS_XOR2X6 U19043 ( .A(w2[5]), .B(n3003), .Z(n8022) );
  HS65_LL_BFX9 U19044 ( .A(n9121), .Z(n9150) );
  HS65_LL_OAI21X3 U19045 ( .A(n3), .B(n1), .C(n2609), .Z(n9111) );
  HS65_LL_IVX9 U19046 ( .A(n2612), .Z(n3) );
  HS65_LL_CBI4I1X5 U19047 ( .A(dcnt[1]), .B(n2610), .C(n2611), .D(dcnt[2]), 
        .Z(n2609) );
  HS65_LL_AO312X9 U19048 ( .A(n5), .B(n4), .C(n2610), .D(n2611), .E(dcnt[1]), 
        .F(n2613), .Z(n9112) );
  HS65_LL_IVX9 U19049 ( .A(dcnt[1]), .Z(n4) );
  HS65_LL_AO22X9 U19050 ( .A(key[109]), .B(n9140), .C(n995), .D(n9149), .Z(
        \u0/N55 ) );
  HS65_LL_AO22X9 U19051 ( .A(key[108]), .B(n9140), .C(n996), .D(n9149), .Z(
        \u0/N54 ) );
  HS65_LL_AO22X9 U19052 ( .A(key[124]), .B(n9141), .C(n980), .D(n9149), .Z(
        \u0/N70 ) );
  HS65_LL_AO22X9 U19053 ( .A(key[100]), .B(n9140), .C(n1004), .D(n9148), .Z(
        \u0/N46 ) );
  HS65_LL_AO22X9 U19054 ( .A(key[116]), .B(n9141), .C(n988), .D(n9143), .Z(
        \u0/N62 ) );
  HS65_LL_AO22X9 U19055 ( .A(key[101]), .B(n9140), .C(n1003), .D(n9143), .Z(
        \u0/N47 ) );
  HS65_LL_AO22X9 U19056 ( .A(key[117]), .B(n9140), .C(n987), .D(n9149), .Z(
        \u0/N63 ) );
endmodule

